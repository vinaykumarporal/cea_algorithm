`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 25.06.2020 09:08:45
// Design Name: 
// Module Name: camellia_F_function
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module camellia_F_function(
    // input are 64-bit FIN and a subkey KE
    input  [63:0] i_fin,
    input  [63:0] i_ke,
    // output is  64-bit FOUT
    output [63:0] o_fout
    );
    
    wire [63:0] w_x;
    
    reg  [7:0] r_t1,
               r_t2,
               r_t3,
               r_t4,
               r_t5,
               r_t6,
               r_t7,
               r_t8;
               
    wire [7:0] w_y1,
               w_y2,
               w_y3,
               w_y4,
               w_y5,
               w_y6,
               w_y7,
               w_y8;
           
    assign w_x = i_fin ^ i_ke;

    always@(*)
        begin
        case(w_x[63:56])
            8'h0   :  r_t1 = 8'h70;
            8'h1   :  r_t1 = 8'h82;
            8'h2   :  r_t1 = 8'h2C;
            8'h3   :  r_t1 = 8'hEC;
            8'h4   :  r_t1 = 8'hB3;
            8'h5   :  r_t1 = 8'h27;
            8'h6   :  r_t1 = 8'hC0;
            8'h7   :  r_t1 = 8'hE5;
            8'h8   :  r_t1 = 8'hE4;
            8'h9   :  r_t1 = 8'h85;
            8'hA   :  r_t1 = 8'h57;
            8'hB   :  r_t1 = 8'h35;
            8'hC   :  r_t1 = 8'hEA;
            8'hD   :  r_t1 = 8'hC;
            8'hE   :  r_t1 = 8'hAE;
            8'hF   :  r_t1 = 8'h41;
            8'h10   :  r_t1 = 8'h23;
            8'h11   :  r_t1 = 8'hEF;
            8'h12   :  r_t1 = 8'h6B;
            8'h13   :  r_t1 = 8'h93;
            8'h14   :  r_t1 = 8'h45;
            8'h15   :  r_t1 = 8'h19;
            8'h16   :  r_t1 = 8'hA5;
            8'h17   :  r_t1 = 8'h21;
            8'h18   :  r_t1 = 8'hED;
            8'h19   :  r_t1 = 8'hE;
            8'h1A   :  r_t1 = 8'h4F;
            8'h1B   :  r_t1 = 8'h4E;
            8'h1C   :  r_t1 = 8'h1D;
            8'h1D   :  r_t1 = 8'h65;
            8'h1E   :  r_t1 = 8'h92;
            8'h1F   :  r_t1 = 8'hBD;
            8'h20   :  r_t1 = 8'h86;
            8'h21   :  r_t1 = 8'hB8;
            8'h22   :  r_t1 = 8'hAF;
            8'h23   :  r_t1 = 8'h8F;
            8'h24   :  r_t1 = 8'h7C;
            8'h25   :  r_t1 = 8'hEB;
            8'h26   :  r_t1 = 8'h1F;
            8'h27   :  r_t1 = 8'hCE;
            8'h28   :  r_t1 = 8'h3E;
            8'h29   :  r_t1 = 8'h30;
            8'h2A   :  r_t1 = 8'hDC;
            8'h2B   :  r_t1 = 8'h5F;
            8'h2C   :  r_t1 = 8'h5E;
            8'h2D   :  r_t1 = 8'hC5;
            8'h2E   :  r_t1 = 8'hB;
            8'h2F   :  r_t1 = 8'h1A;
            8'h30   :  r_t1 = 8'hA6;
            8'h31   :  r_t1 = 8'hE1;
            8'h32   :  r_t1 = 8'h39;
            8'h33   :  r_t1 = 8'hCA;
            8'h34   :  r_t1 = 8'hD5;
            8'h35   :  r_t1 = 8'h47;
            8'h36   :  r_t1 = 8'h5D;
            8'h37   :  r_t1 = 8'h3D;
            8'h38   :  r_t1 = 8'hD9;
            8'h39   :  r_t1 = 8'h1;
            8'h3A   :  r_t1 = 8'h5A;
            8'h3B   :  r_t1 = 8'hD6;
            8'h3C   :  r_t1 = 8'h51;
            8'h3D   :  r_t1 = 8'h56;
            8'h3E   :  r_t1 = 8'h6C;
            8'h3F   :  r_t1 = 8'h4D;
            8'h40   :  r_t1 = 8'h8B;
            8'h41   :  r_t1 = 8'hD;
            8'h42   :  r_t1 = 8'h9A;
            8'h43   :  r_t1 = 8'h66;
            8'h44   :  r_t1 = 8'hFB;
            8'h45   :  r_t1 = 8'hCC;
            8'h46   :  r_t1 = 8'hB0;
            8'h47   :  r_t1 = 8'h2D;
            8'h48   :  r_t1 = 8'h74;
            8'h49   :  r_t1 = 8'h12;
            8'h4A   :  r_t1 = 8'h2B;
            8'h4B   :  r_t1 = 8'h20;
            8'h4C   :  r_t1 = 8'hF0;
            8'h4D   :  r_t1 = 8'hB1;
            8'h4E   :  r_t1 = 8'h84;
            8'h4F   :  r_t1 = 8'h99;
            8'h50   :  r_t1 = 8'hDF;
            8'h51   :  r_t1 = 8'h4C;
            8'h52   :  r_t1 = 8'hCB;
            8'h53   :  r_t1 = 8'hC2;
            8'h54   :  r_t1 = 8'h34;
            8'h55   :  r_t1 = 8'h7E;
            8'h56   :  r_t1 = 8'h76;
            8'h57   :  r_t1 = 8'h5;
            8'h58   :  r_t1 = 8'h6D;
            8'h59   :  r_t1 = 8'hB7;
            8'h5A   :  r_t1 = 8'hA9;
            8'h5B   :  r_t1 = 8'h31;
            8'h5C   :  r_t1 = 8'hD1;
            8'h5D   :  r_t1 = 8'h17;
            8'h5E   :  r_t1 = 8'h4;
            8'h5F   :  r_t1 = 8'hD7;
            8'h60   :  r_t1 = 8'h14;
            8'h61   :  r_t1 = 8'h58;
            8'h62   :  r_t1 = 8'h3A;
            8'h63   :  r_t1 = 8'h61;
            8'h64   :  r_t1 = 8'hDE;
            8'h65   :  r_t1 = 8'h1B;
            8'h66   :  r_t1 = 8'h11;
            8'h67   :  r_t1 = 8'h1C;
            8'h68   :  r_t1 = 8'h32;
            8'h69   :  r_t1 = 8'hF;
            8'h6A   :  r_t1 = 8'h9C;
            8'h6B   :  r_t1 = 8'h16;
            8'h6C   :  r_t1 = 8'h53;
            8'h6D   :  r_t1 = 8'h18;
            8'h6E   :  r_t1 = 8'hF2;
            8'h6F   :  r_t1 = 8'h22;
            8'h70   :  r_t1 = 8'hFE;
            8'h71   :  r_t1 = 8'h44;
            8'h72   :  r_t1 = 8'hCF;
            8'h73   :  r_t1 = 8'hB2;
            8'h74   :  r_t1 = 8'hC3;
            8'h75   :  r_t1 = 8'hB5;
            8'h76   :  r_t1 = 8'h7A;
            8'h77   :  r_t1 = 8'h91;
            8'h78   :  r_t1 = 8'h24;
            8'h79   :  r_t1 = 8'h8;
            8'h7A   :  r_t1 = 8'hE8;
            8'h7B   :  r_t1 = 8'hA8;
            8'h7C   :  r_t1 = 8'h60;
            8'h7D   :  r_t1 = 8'hFC;
            8'h7E   :  r_t1 = 8'h69;
            8'h7F   :  r_t1 = 8'h50;
            8'h80   :  r_t1 = 8'hAA;
            8'h81   :  r_t1 = 8'hD0;
            8'h82   :  r_t1 = 8'hA0;
            8'h83   :  r_t1 = 8'h7D;
            8'h84   :  r_t1 = 8'hA1;
            8'h85   :  r_t1 = 8'h89;
            8'h86   :  r_t1 = 8'h62;
            8'h87   :  r_t1 = 8'h97;
            8'h88   :  r_t1 = 8'h54;
            8'h89   :  r_t1 = 8'h5B;
            8'h8A   :  r_t1 = 8'h1E;
            8'h8B   :  r_t1 = 8'h95;
            8'h8C   :  r_t1 = 8'hE0;
            8'h8D   :  r_t1 = 8'hFF;
            8'h8E   :  r_t1 = 8'h64;
            8'h8F   :  r_t1 = 8'hD2;
            8'h90   :  r_t1 = 8'h10;
            8'h91   :  r_t1 = 8'hC4;
            8'h92   :  r_t1 = 8'h0;
            8'h93   :  r_t1 = 8'h48;
            8'h94   :  r_t1 = 8'hA3;
            8'h95   :  r_t1 = 8'hF7;
            8'h96   :  r_t1 = 8'h75;
            8'h97   :  r_t1 = 8'hDB;
            8'h98   :  r_t1 = 8'h8A;
            8'h99   :  r_t1 = 8'h3;
            8'h9A   :  r_t1 = 8'hE6;
            8'h9B   :  r_t1 = 8'hDA;
            8'h9C   :  r_t1 = 8'h9;
            8'h9D   :  r_t1 = 8'h3F;
            8'h9E   :  r_t1 = 8'hDD;
            8'h9F   :  r_t1 = 8'h94;
            8'hA0   :  r_t1 = 8'h87;
            8'hA1   :  r_t1 = 8'h5C;
            8'hA2   :  r_t1 = 8'h83;
            8'hA3   :  r_t1 = 8'h2;
            8'hA4   :  r_t1 = 8'hCD;
            8'hA5   :  r_t1 = 8'h4A;
            8'hA6   :  r_t1 = 8'h90;
            8'hA7   :  r_t1 = 8'h33;
            8'hA8   :  r_t1 = 8'h73;
            8'hA9   :  r_t1 = 8'h67;
            8'hAA   :  r_t1 = 8'hF6;
            8'hAB   :  r_t1 = 8'hF3;
            8'hAC   :  r_t1 = 8'h9D;
            8'hAD   :  r_t1 = 8'h7F;
            8'hAE   :  r_t1 = 8'hBF;
            8'hAF   :  r_t1 = 8'hE2;
            8'hB0   :  r_t1 = 8'h52;
            8'hB1   :  r_t1 = 8'h9B;
            8'hB2   :  r_t1 = 8'hD8;
            8'hB3   :  r_t1 = 8'h26;
            8'hB4   :  r_t1 = 8'hC8;
            8'hB5   :  r_t1 = 8'h37;
            8'hB6   :  r_t1 = 8'hC6;
            8'hB7   :  r_t1 = 8'h3B;
            8'hB8   :  r_t1 = 8'h81;
            8'hB9   :  r_t1 = 8'h96;
            8'hBA   :  r_t1 = 8'h6F;
            8'hBB   :  r_t1 = 8'h4B;
            8'hBC   :  r_t1 = 8'h13;
            8'hBD   :  r_t1 = 8'hBE;
            8'hBE   :  r_t1 = 8'h63;
            8'hBF   :  r_t1 = 8'h2E;
            8'hC0   :  r_t1 = 8'hE9;
            8'hC1   :  r_t1 = 8'h79;
            8'hC2   :  r_t1 = 8'hA7;
            8'hC3   :  r_t1 = 8'h8C;
            8'hC4   :  r_t1 = 8'h9F;
            8'hC5   :  r_t1 = 8'h6E;
            8'hC6   :  r_t1 = 8'hBC;
            8'hC7   :  r_t1 = 8'h8E;
            8'hC8   :  r_t1 = 8'h29;
            8'hC9   :  r_t1 = 8'hF5;
            8'hCA   :  r_t1 = 8'hF9;
            8'hCB   :  r_t1 = 8'hB6;
            8'hCC   :  r_t1 = 8'h2F;
            8'hCD   :  r_t1 = 8'hFD;
            8'hCE   :  r_t1 = 8'hB4;
            8'hCF   :  r_t1 = 8'h59;
            8'hD0   :  r_t1 = 8'h78;
            8'hD1   :  r_t1 = 8'h98;
            8'hD2   :  r_t1 = 8'h6;
            8'hD3   :  r_t1 = 8'h6A;
            8'hD4   :  r_t1 = 8'hE7;
            8'hD5   :  r_t1 = 8'h46;
            8'hD6   :  r_t1 = 8'h71;
            8'hD7   :  r_t1 = 8'hBA;
            8'hD8   :  r_t1 = 8'hD4;
            8'hD9   :  r_t1 = 8'h25;
            8'hDA   :  r_t1 = 8'hAB;
            8'hDB   :  r_t1 = 8'h42;
            8'hDC   :  r_t1 = 8'h88;
            8'hDD   :  r_t1 = 8'hA2;
            8'hDE   :  r_t1 = 8'h8D;
            8'hDF   :  r_t1 = 8'hFA;
            8'hE0   :  r_t1 = 8'h72;
            8'hE1   :  r_t1 = 8'h7;
            8'hE2   :  r_t1 = 8'hB9;
            8'hE3   :  r_t1 = 8'h55;
            8'hE4   :  r_t1 = 8'hF8;
            8'hE5   :  r_t1 = 8'hEE;
            8'hE6   :  r_t1 = 8'hAC;
            8'hE7   :  r_t1 = 8'hA;
            8'hE8   :  r_t1 = 8'h36;
            8'hE9   :  r_t1 = 8'h49;
            8'hEA   :  r_t1 = 8'h2A;
            8'hEB   :  r_t1 = 8'h68;
            8'hEC   :  r_t1 = 8'h3C;
            8'hED   :  r_t1 = 8'h38;
            8'hEE   :  r_t1 = 8'hF1;
            8'hEF   :  r_t1 = 8'hA4;
            8'hF0   :  r_t1 = 8'h40;
            8'hF1   :  r_t1 = 8'h28;
            8'hF2   :  r_t1 = 8'hD3;
            8'hF3   :  r_t1 = 8'h7B;
            8'hF4   :  r_t1 = 8'hBB;
            8'hF5   :  r_t1 = 8'hC9;
            8'hF6   :  r_t1 = 8'h43;
            8'hF7   :  r_t1 = 8'hC1;
            8'hF8   :  r_t1 = 8'h15;
            8'hF9   :  r_t1 = 8'hE3;
            8'hFA   :  r_t1 = 8'hAD;
            8'hFB   :  r_t1 = 8'hF4;
            8'hFC   :  r_t1 = 8'h77;
            8'hFD   :  r_t1 = 8'hC7;
            8'hFE   :  r_t1 = 8'h80;
            8'hFF   :  r_t1 = 8'h9E;
        endcase
        end
        
    always@(*)
        begin
        case(w_x[55:48])
            8'h0   :  r_t2 = 8'hE0;
            8'h1   :  r_t2 = 8'h5;
            8'h2   :  r_t2 = 8'h58;
            8'h3   :  r_t2 = 8'hD9;
            8'h4   :  r_t2 = 8'h67;
            8'h5   :  r_t2 = 8'h4E;
            8'h6   :  r_t2 = 8'h81;
            8'h7   :  r_t2 = 8'hCB;
            8'h8   :  r_t2 = 8'hC9;
            8'h9   :  r_t2 = 8'hB;
            8'hA   :  r_t2 = 8'hAE;
            8'hB   :  r_t2 = 8'h6A;
            8'hC   :  r_t2 = 8'hD5;
            8'hD   :  r_t2 = 8'h18;
            8'hE   :  r_t2 = 8'h5D;
            8'hF   :  r_t2 = 8'h82;
            8'h10   :  r_t2 = 8'h46;
            8'h11   :  r_t2 = 8'hDF;
            8'h12   :  r_t2 = 8'hD6;
            8'h13   :  r_t2 = 8'h27;
            8'h14   :  r_t2 = 8'h8A;
            8'h15   :  r_t2 = 8'h32;
            8'h16   :  r_t2 = 8'h4B;
            8'h17   :  r_t2 = 8'h42;
            8'h18   :  r_t2 = 8'hDB;
            8'h19   :  r_t2 = 8'h1C;
            8'h1A   :  r_t2 = 8'h9E;
            8'h1B   :  r_t2 = 8'h9C;
            8'h1C   :  r_t2 = 8'h3A;
            8'h1D   :  r_t2 = 8'hCA;
            8'h1E   :  r_t2 = 8'h25;
            8'h1F   :  r_t2 = 8'h7B;
            8'h20   :  r_t2 = 8'hD;
            8'h21   :  r_t2 = 8'h71;
            8'h22   :  r_t2 = 8'h5F;
            8'h23   :  r_t2 = 8'h1F;
            8'h24   :  r_t2 = 8'hF8;
            8'h25   :  r_t2 = 8'hD7;
            8'h26   :  r_t2 = 8'h3E;
            8'h27   :  r_t2 = 8'h9D;
            8'h28   :  r_t2 = 8'h7C;
            8'h29   :  r_t2 = 8'h60;
            8'h2A   :  r_t2 = 8'hB9;
            8'h2B   :  r_t2 = 8'hBE;
            8'h2C   :  r_t2 = 8'hBC;
            8'h2D   :  r_t2 = 8'h8B;
            8'h2E   :  r_t2 = 8'h16;
            8'h2F   :  r_t2 = 8'h34;
            8'h30   :  r_t2 = 8'h4D;
            8'h31   :  r_t2 = 8'hC3;
            8'h32   :  r_t2 = 8'h72;
            8'h33   :  r_t2 = 8'h95;
            8'h34   :  r_t2 = 8'hAB;
            8'h35   :  r_t2 = 8'h8E;
            8'h36   :  r_t2 = 8'hBA;
            8'h37   :  r_t2 = 8'h7A;
            8'h38   :  r_t2 = 8'hB3;
            8'h39   :  r_t2 = 8'h2;
            8'h3A   :  r_t2 = 8'hB4;
            8'h3B   :  r_t2 = 8'hAD;
            8'h3C   :  r_t2 = 8'hA2;
            8'h3D   :  r_t2 = 8'hAC;
            8'h3E   :  r_t2 = 8'hD8;
            8'h3F   :  r_t2 = 8'h9A;
            8'h40   :  r_t2 = 8'h17;
            8'h41   :  r_t2 = 8'h1A;
            8'h42   :  r_t2 = 8'h35;
            8'h43   :  r_t2 = 8'hCC;
            8'h44   :  r_t2 = 8'hF7;
            8'h45   :  r_t2 = 8'h99;
            8'h46   :  r_t2 = 8'h61;
            8'h47   :  r_t2 = 8'h5A;
            8'h48   :  r_t2 = 8'hE8;
            8'h49   :  r_t2 = 8'h24;
            8'h4A   :  r_t2 = 8'h56;
            8'h4B   :  r_t2 = 8'h40;
            8'h4C   :  r_t2 = 8'hE1;
            8'h4D   :  r_t2 = 8'h63;
            8'h4E   :  r_t2 = 8'h9;
            8'h4F   :  r_t2 = 8'h33;
            8'h50   :  r_t2 = 8'hBF;
            8'h51   :  r_t2 = 8'h98;
            8'h52   :  r_t2 = 8'h97;
            8'h53   :  r_t2 = 8'h85;
            8'h54   :  r_t2 = 8'h68;
            8'h55   :  r_t2 = 8'hFC;
            8'h56   :  r_t2 = 8'hEC;
            8'h57   :  r_t2 = 8'hA;
            8'h58   :  r_t2 = 8'hDA;
            8'h59   :  r_t2 = 8'h6F;
            8'h5A   :  r_t2 = 8'h53;
            8'h5B   :  r_t2 = 8'h62;
            8'h5C   :  r_t2 = 8'hA3;
            8'h5D   :  r_t2 = 8'h2E;
            8'h5E   :  r_t2 = 8'h8;
            8'h5F   :  r_t2 = 8'hAF;
            8'h60   :  r_t2 = 8'h28;
            8'h61   :  r_t2 = 8'hB0;
            8'h62   :  r_t2 = 8'h74;
            8'h63   :  r_t2 = 8'hC2;
            8'h64   :  r_t2 = 8'hBD;
            8'h65   :  r_t2 = 8'h36;
            8'h66   :  r_t2 = 8'h22;
            8'h67   :  r_t2 = 8'h38;
            8'h68   :  r_t2 = 8'h64;
            8'h69   :  r_t2 = 8'h1E;
            8'h6A   :  r_t2 = 8'h39;
            8'h6B   :  r_t2 = 8'h2C;
            8'h6C   :  r_t2 = 8'hA6;
            8'h6D   :  r_t2 = 8'h30;
            8'h6E   :  r_t2 = 8'hE5;
            8'h6F   :  r_t2 = 8'h44;
            8'h70   :  r_t2 = 8'hFD;
            8'h71   :  r_t2 = 8'h88;
            8'h72   :  r_t2 = 8'h9F;
            8'h73   :  r_t2 = 8'h65;
            8'h74   :  r_t2 = 8'h87;
            8'h75   :  r_t2 = 8'h6B;
            8'h76   :  r_t2 = 8'hF4;
            8'h77   :  r_t2 = 8'h23;
            8'h78   :  r_t2 = 8'h48;
            8'h79   :  r_t2 = 8'h10;
            8'h7A   :  r_t2 = 8'hD1;
            8'h7B   :  r_t2 = 8'h51;
            8'h7C   :  r_t2 = 8'hC0;
            8'h7D   :  r_t2 = 8'hF9;
            8'h7E   :  r_t2 = 8'hD2;
            8'h7F   :  r_t2 = 8'hA0;
            8'h80   :  r_t2 = 8'h55;
            8'h81   :  r_t2 = 8'hA1;
            8'h82   :  r_t2 = 8'h41;
            8'h83   :  r_t2 = 8'hFA;
            8'h84   :  r_t2 = 8'h43;
            8'h85   :  r_t2 = 8'h13;
            8'h86   :  r_t2 = 8'hC4;
            8'h87   :  r_t2 = 8'h2F;
            8'h88   :  r_t2 = 8'hA8;
            8'h89   :  r_t2 = 8'hB6;
            8'h8A   :  r_t2 = 8'h3C;
            8'h8B   :  r_t2 = 8'h2B;
            8'h8C   :  r_t2 = 8'hC1;
            8'h8D   :  r_t2 = 8'hFF;
            8'h8E   :  r_t2 = 8'hC8;
            8'h8F   :  r_t2 = 8'hA5;
            8'h90   :  r_t2 = 8'h20;
            8'h91   :  r_t2 = 8'h89;
            8'h92   :  r_t2 = 8'h0;
            8'h93   :  r_t2 = 8'h90;
            8'h94   :  r_t2 = 8'h47;
            8'h95   :  r_t2 = 8'hEF;
            8'h96   :  r_t2 = 8'hEA;
            8'h97   :  r_t2 = 8'hB7;
            8'h98   :  r_t2 = 8'h15;
            8'h99   :  r_t2 = 8'h6;
            8'h9A   :  r_t2 = 8'hCD;
            8'h9B   :  r_t2 = 8'hB5;
            8'h9C   :  r_t2 = 8'h12;
            8'h9D   :  r_t2 = 8'h7E;
            8'h9E   :  r_t2 = 8'hBB;
            8'h9F   :  r_t2 = 8'h29;
            8'hA0   :  r_t2 = 8'hF;
            8'hA1   :  r_t2 = 8'hB8;
            8'hA2   :  r_t2 = 8'h7;
            8'hA3   :  r_t2 = 8'h4;
            8'hA4   :  r_t2 = 8'h9B;
            8'hA5   :  r_t2 = 8'h94;
            8'hA6   :  r_t2 = 8'h21;
            8'hA7   :  r_t2 = 8'h66;
            8'hA8   :  r_t2 = 8'hE6;
            8'hA9   :  r_t2 = 8'hCE;
            8'hAA   :  r_t2 = 8'hED;
            8'hAB   :  r_t2 = 8'hE7;
            8'hAC   :  r_t2 = 8'h3B;
            8'hAD   :  r_t2 = 8'hFE;
            8'hAE   :  r_t2 = 8'h7F;
            8'hAF   :  r_t2 = 8'hC5;
            8'hB0   :  r_t2 = 8'hA4;
            8'hB1   :  r_t2 = 8'h37;
            8'hB2   :  r_t2 = 8'hB1;
            8'hB3   :  r_t2 = 8'h4C;
            8'hB4   :  r_t2 = 8'h91;
            8'hB5   :  r_t2 = 8'h6E;
            8'hB6   :  r_t2 = 8'h8D;
            8'hB7   :  r_t2 = 8'h76;
            8'hB8   :  r_t2 = 8'h3;
            8'hB9   :  r_t2 = 8'h2D;
            8'hBA   :  r_t2 = 8'hDE;
            8'hBB   :  r_t2 = 8'h96;
            8'hBC   :  r_t2 = 8'h26;
            8'hBD   :  r_t2 = 8'h7D;
            8'hBE   :  r_t2 = 8'hC6;
            8'hBF   :  r_t2 = 8'h5C;
            8'hC0   :  r_t2 = 8'hD3;
            8'hC1   :  r_t2 = 8'hF2;
            8'hC2   :  r_t2 = 8'h4F;
            8'hC3   :  r_t2 = 8'h19;
            8'hC4   :  r_t2 = 8'h3F;
            8'hC5   :  r_t2 = 8'hDC;
            8'hC6   :  r_t2 = 8'h79;
            8'hC7   :  r_t2 = 8'h1D;
            8'hC8   :  r_t2 = 8'h52;
            8'hC9   :  r_t2 = 8'hEB;
            8'hCA   :  r_t2 = 8'hF3;
            8'hCB   :  r_t2 = 8'h6D;
            8'hCC   :  r_t2 = 8'h5E;
            8'hCD   :  r_t2 = 8'hFB;
            8'hCE   :  r_t2 = 8'h69;
            8'hCF   :  r_t2 = 8'hB2;
            8'hD0   :  r_t2 = 8'hF0;
            8'hD1   :  r_t2 = 8'h31;
            8'hD2   :  r_t2 = 8'hC;
            8'hD3   :  r_t2 = 8'hD4;
            8'hD4   :  r_t2 = 8'hCF;
            8'hD5   :  r_t2 = 8'h8C;
            8'hD6   :  r_t2 = 8'hE2;
            8'hD7   :  r_t2 = 8'h75;
            8'hD8   :  r_t2 = 8'hA9;
            8'hD9   :  r_t2 = 8'h4A;
            8'hDA   :  r_t2 = 8'h57;
            8'hDB   :  r_t2 = 8'h84;
            8'hDC   :  r_t2 = 8'h11;
            8'hDD   :  r_t2 = 8'h45;
            8'hDE   :  r_t2 = 8'h1B;
            8'hDF   :  r_t2 = 8'hF5;
            8'hE0   :  r_t2 = 8'hE4;
            8'hE1   :  r_t2 = 8'hE;
            8'hE2   :  r_t2 = 8'h73;
            8'hE3   :  r_t2 = 8'hAA;
            8'hE4   :  r_t2 = 8'hF1;
            8'hE5   :  r_t2 = 8'hDD;
            8'hE6   :  r_t2 = 8'h59;
            8'hE7   :  r_t2 = 8'h14;
            8'hE8   :  r_t2 = 8'h6C;
            8'hE9   :  r_t2 = 8'h92;
            8'hEA   :  r_t2 = 8'h54;
            8'hEB   :  r_t2 = 8'hD0;
            8'hEC   :  r_t2 = 8'h78;
            8'hED   :  r_t2 = 8'h70;
            8'hEE   :  r_t2 = 8'hE3;
            8'hEF   :  r_t2 = 8'h49;
            8'hF0   :  r_t2 = 8'h80;
            8'hF1   :  r_t2 = 8'h50;
            8'hF2   :  r_t2 = 8'hA7;
            8'hF3   :  r_t2 = 8'hF6;
            8'hF4   :  r_t2 = 8'h77;
            8'hF5   :  r_t2 = 8'h93;
            8'hF6   :  r_t2 = 8'h86;
            8'hF7   :  r_t2 = 8'h83;
            8'hF8   :  r_t2 = 8'h2A;
            8'hF9   :  r_t2 = 8'hC7;
            8'hFA   :  r_t2 = 8'h5B;
            8'hFB   :  r_t2 = 8'hE9;
            8'hFC   :  r_t2 = 8'hEE;
            8'hFD   :  r_t2 = 8'h8F;
            8'hFE   :  r_t2 = 8'h1;
            8'hFF   :  r_t2 = 8'h3D;
        endcase
        end
        
    always@(*)
        begin
        case(w_x[47:40])
            8'h0   :  r_t3 = 8'h38;
            8'h1   :  r_t3 = 8'h41;
            8'h2   :  r_t3 = 8'h16;
            8'h3   :  r_t3 = 8'h76;
            8'h4   :  r_t3 = 8'hD9;
            8'h5   :  r_t3 = 8'h93;
            8'h6   :  r_t3 = 8'h60;
            8'h7   :  r_t3 = 8'hF2;
            8'h8   :  r_t3 = 8'h72;
            8'h9   :  r_t3 = 8'hC2;
            8'hA   :  r_t3 = 8'hAB;
            8'hB   :  r_t3 = 8'h9A;
            8'hC   :  r_t3 = 8'h75;
            8'hD   :  r_t3 = 8'h6;
            8'hE   :  r_t3 = 8'h57;
            8'hF   :  r_t3 = 8'hA0;
            8'h10   :  r_t3 = 8'h91;
            8'h11   :  r_t3 = 8'hF7;
            8'h12   :  r_t3 = 8'hB5;
            8'h13   :  r_t3 = 8'hC9;
            8'h14   :  r_t3 = 8'hA2;
            8'h15   :  r_t3 = 8'h8C;
            8'h16   :  r_t3 = 8'hD2;
            8'h17   :  r_t3 = 8'h90;
            8'h18   :  r_t3 = 8'hF6;
            8'h19   :  r_t3 = 8'h7;
            8'h1A   :  r_t3 = 8'hA7;
            8'h1B   :  r_t3 = 8'h27;
            8'h1C   :  r_t3 = 8'h8E;
            8'h1D   :  r_t3 = 8'hB2;
            8'h1E   :  r_t3 = 8'h49;
            8'h1F   :  r_t3 = 8'hDE;
            8'h20   :  r_t3 = 8'h43;
            8'h21   :  r_t3 = 8'h5C;
            8'h22   :  r_t3 = 8'hD7;
            8'h23   :  r_t3 = 8'hC7;
            8'h24   :  r_t3 = 8'h3E;
            8'h25   :  r_t3 = 8'hF5;
            8'h26   :  r_t3 = 8'h8F;
            8'h27   :  r_t3 = 8'h67;
            8'h28   :  r_t3 = 8'h1F;
            8'h29   :  r_t3 = 8'h18;
            8'h2A   :  r_t3 = 8'h6E;
            8'h2B   :  r_t3 = 8'hAF;
            8'h2C   :  r_t3 = 8'h2F;
            8'h2D   :  r_t3 = 8'hE2;
            8'h2E   :  r_t3 = 8'h85;
            8'h2F   :  r_t3 = 8'hD;
            8'h30   :  r_t3 = 8'h53;
            8'h31   :  r_t3 = 8'hF0;
            8'h32   :  r_t3 = 8'h9C;
            8'h33   :  r_t3 = 8'h65;
            8'h34   :  r_t3 = 8'hEA;
            8'h35   :  r_t3 = 8'hA3;
            8'h36   :  r_t3 = 8'hAE;
            8'h37   :  r_t3 = 8'h9E;
            8'h38   :  r_t3 = 8'hEC;
            8'h39   :  r_t3 = 8'h80;
            8'h3A   :  r_t3 = 8'h2D;
            8'h3B   :  r_t3 = 8'h6B;
            8'h3C   :  r_t3 = 8'hA8;
            8'h3D   :  r_t3 = 8'h2B;
            8'h3E   :  r_t3 = 8'h36;
            8'h3F   :  r_t3 = 8'hA6;
            8'h40   :  r_t3 = 8'hC5;
            8'h41   :  r_t3 = 8'h86;
            8'h42   :  r_t3 = 8'h4D;
            8'h43   :  r_t3 = 8'h33;
            8'h44   :  r_t3 = 8'hFD;
            8'h45   :  r_t3 = 8'h66;
            8'h46   :  r_t3 = 8'h58;
            8'h47   :  r_t3 = 8'h96;
            8'h48   :  r_t3 = 8'h3A;
            8'h49   :  r_t3 = 8'h9;
            8'h4A   :  r_t3 = 8'h95;
            8'h4B   :  r_t3 = 8'h10;
            8'h4C   :  r_t3 = 8'h78;
            8'h4D   :  r_t3 = 8'hD8;
            8'h4E   :  r_t3 = 8'h42;
            8'h4F   :  r_t3 = 8'hCC;
            8'h50   :  r_t3 = 8'hEF;
            8'h51   :  r_t3 = 8'h26;
            8'h52   :  r_t3 = 8'hE5;
            8'h53   :  r_t3 = 8'h61;
            8'h54   :  r_t3 = 8'h1A;
            8'h55   :  r_t3 = 8'h3F;
            8'h56   :  r_t3 = 8'h3B;
            8'h57   :  r_t3 = 8'h82;
            8'h58   :  r_t3 = 8'hB6;
            8'h59   :  r_t3 = 8'hDB;
            8'h5A   :  r_t3 = 8'hD4;
            8'h5B   :  r_t3 = 8'h98;
            8'h5C   :  r_t3 = 8'hE8;
            8'h5D   :  r_t3 = 8'h8B;
            8'h5E   :  r_t3 = 8'h2;
            8'h5F   :  r_t3 = 8'hEB;
            8'h60   :  r_t3 = 8'hA;
            8'h61   :  r_t3 = 8'h2C;
            8'h62   :  r_t3 = 8'h1D;
            8'h63   :  r_t3 = 8'hB0;
            8'h64   :  r_t3 = 8'h6F;
            8'h65   :  r_t3 = 8'h8D;
            8'h66   :  r_t3 = 8'h88;
            8'h67   :  r_t3 = 8'hE;
            8'h68   :  r_t3 = 8'h19;
            8'h69   :  r_t3 = 8'h87;
            8'h6A   :  r_t3 = 8'h4E;
            8'h6B   :  r_t3 = 8'hB;
            8'h6C   :  r_t3 = 8'hA9;
            8'h6D   :  r_t3 = 8'hC;
            8'h6E   :  r_t3 = 8'h79;
            8'h6F   :  r_t3 = 8'h11;
            8'h70   :  r_t3 = 8'h7F;
            8'h71   :  r_t3 = 8'h22;
            8'h72   :  r_t3 = 8'hE7;
            8'h73   :  r_t3 = 8'h59;
            8'h74   :  r_t3 = 8'hE1;
            8'h75   :  r_t3 = 8'hDA;
            8'h76   :  r_t3 = 8'h3D;
            8'h77   :  r_t3 = 8'hC8;
            8'h78   :  r_t3 = 8'h12;
            8'h79   :  r_t3 = 8'h4;
            8'h7A   :  r_t3 = 8'h74;
            8'h7B   :  r_t3 = 8'h54;
            8'h7C   :  r_t3 = 8'h30;
            8'h7D   :  r_t3 = 8'h7E;
            8'h7E   :  r_t3 = 8'hB4;
            8'h7F   :  r_t3 = 8'h28;
            8'h80   :  r_t3 = 8'h55;
            8'h81   :  r_t3 = 8'h68;
            8'h82   :  r_t3 = 8'h50;
            8'h83   :  r_t3 = 8'hBE;
            8'h84   :  r_t3 = 8'hD0;
            8'h85   :  r_t3 = 8'hC4;
            8'h86   :  r_t3 = 8'h31;
            8'h87   :  r_t3 = 8'hCB;
            8'h88   :  r_t3 = 8'h2A;
            8'h89   :  r_t3 = 8'hAD;
            8'h8A   :  r_t3 = 8'hF;
            8'h8B   :  r_t3 = 8'hCA;
            8'h8C   :  r_t3 = 8'h70;
            8'h8D   :  r_t3 = 8'hFF;
            8'h8E   :  r_t3 = 8'h32;
            8'h8F   :  r_t3 = 8'h69;
            8'h90   :  r_t3 = 8'h8;
            8'h91   :  r_t3 = 8'h62;
            8'h92   :  r_t3 = 8'h0;
            8'h93   :  r_t3 = 8'h24;
            8'h94   :  r_t3 = 8'hD1;
            8'h95   :  r_t3 = 8'hFB;
            8'h96   :  r_t3 = 8'hBA;
            8'h97   :  r_t3 = 8'hED;
            8'h98   :  r_t3 = 8'h45;
            8'h99   :  r_t3 = 8'h81;
            8'h9A   :  r_t3 = 8'h73;
            8'h9B   :  r_t3 = 8'h6D;
            8'h9C   :  r_t3 = 8'h84;
            8'h9D   :  r_t3 = 8'h9F;
            8'h9E   :  r_t3 = 8'hEE;
            8'h9F   :  r_t3 = 8'h4A;
            8'hA0   :  r_t3 = 8'hC3;
            8'hA1   :  r_t3 = 8'h2E;
            8'hA2   :  r_t3 = 8'hC1;
            8'hA3   :  r_t3 = 8'h1;
            8'hA4   :  r_t3 = 8'hE6;
            8'hA5   :  r_t3 = 8'h25;
            8'hA6   :  r_t3 = 8'h48;
            8'hA7   :  r_t3 = 8'h99;
            8'hA8   :  r_t3 = 8'hB9;
            8'hA9   :  r_t3 = 8'hB3;
            8'hAA   :  r_t3 = 8'h7B;
            8'hAB   :  r_t3 = 8'hF9;
            8'hAC   :  r_t3 = 8'hCE;
            8'hAD   :  r_t3 = 8'hBF;
            8'hAE   :  r_t3 = 8'hDF;
            8'hAF   :  r_t3 = 8'h71;
            8'hB0   :  r_t3 = 8'h29;
            8'hB1   :  r_t3 = 8'hCD;
            8'hB2   :  r_t3 = 8'h6C;
            8'hB3   :  r_t3 = 8'h13;
            8'hB4   :  r_t3 = 8'h64;
            8'hB5   :  r_t3 = 8'h9B;
            8'hB6   :  r_t3 = 8'h63;
            8'hB7   :  r_t3 = 8'h9D;
            8'hB8   :  r_t3 = 8'hC0;
            8'hB9   :  r_t3 = 8'h4B;
            8'hBA   :  r_t3 = 8'hB7;
            8'hBB   :  r_t3 = 8'hA5;
            8'hBC   :  r_t3 = 8'h89;
            8'hBD   :  r_t3 = 8'h5F;
            8'hBE   :  r_t3 = 8'hB1;
            8'hBF   :  r_t3 = 8'h17;
            8'hC0   :  r_t3 = 8'hF4;
            8'hC1   :  r_t3 = 8'hBC;
            8'hC2   :  r_t3 = 8'hD3;
            8'hC3   :  r_t3 = 8'h46;
            8'hC4   :  r_t3 = 8'hCF;
            8'hC5   :  r_t3 = 8'h37;
            8'hC6   :  r_t3 = 8'h5E;
            8'hC7   :  r_t3 = 8'h47;
            8'hC8   :  r_t3 = 8'h94;
            8'hC9   :  r_t3 = 8'hFA;
            8'hCA   :  r_t3 = 8'hFC;
            8'hCB   :  r_t3 = 8'h5B;
            8'hCC   :  r_t3 = 8'h97;
            8'hCD   :  r_t3 = 8'hFE;
            8'hCE   :  r_t3 = 8'h5A;
            8'hCF   :  r_t3 = 8'hAC;
            8'hD0   :  r_t3 = 8'h3C;
            8'hD1   :  r_t3 = 8'h4C;
            8'hD2   :  r_t3 = 8'h3;
            8'hD3   :  r_t3 = 8'h35;
            8'hD4   :  r_t3 = 8'hF3;
            8'hD5   :  r_t3 = 8'h23;
            8'hD6   :  r_t3 = 8'hB8;
            8'hD7   :  r_t3 = 8'h5D;
            8'hD8   :  r_t3 = 8'h6A;
            8'hD9   :  r_t3 = 8'h92;
            8'hDA   :  r_t3 = 8'hD5;
            8'hDB   :  r_t3 = 8'h21;
            8'hDC   :  r_t3 = 8'h44;
            8'hDD   :  r_t3 = 8'h51;
            8'hDE   :  r_t3 = 8'hC6;
            8'hDF   :  r_t3 = 8'h7D;
            8'hE0   :  r_t3 = 8'h39;
            8'hE1   :  r_t3 = 8'h83;
            8'hE2   :  r_t3 = 8'hDC;
            8'hE3   :  r_t3 = 8'hAA;
            8'hE4   :  r_t3 = 8'h7C;
            8'hE5   :  r_t3 = 8'h77;
            8'hE6   :  r_t3 = 8'h56;
            8'hE7   :  r_t3 = 8'h5;
            8'hE8   :  r_t3 = 8'h1B;
            8'hE9   :  r_t3 = 8'hA4;
            8'hEA   :  r_t3 = 8'h15;
            8'hEB   :  r_t3 = 8'h34;
            8'hEC   :  r_t3 = 8'h1E;
            8'hED   :  r_t3 = 8'h1C;
            8'hEE   :  r_t3 = 8'hF8;
            8'hEF   :  r_t3 = 8'h52;
            8'hF0   :  r_t3 = 8'h20;
            8'hF1   :  r_t3 = 8'h14;
            8'hF2   :  r_t3 = 8'hE9;
            8'hF3   :  r_t3 = 8'hBD;
            8'hF4   :  r_t3 = 8'hDD;
            8'hF5   :  r_t3 = 8'hE4;
            8'hF6   :  r_t3 = 8'hA1;
            8'hF7   :  r_t3 = 8'hE0;
            8'hF8   :  r_t3 = 8'h8A;
            8'hF9   :  r_t3 = 8'hF1;
            8'hFA   :  r_t3 = 8'hD6;
            8'hFB   :  r_t3 = 8'h7A;
            8'hFC   :  r_t3 = 8'hBB;
            8'hFD   :  r_t3 = 8'hE3;
            8'hFE   :  r_t3 = 8'h40;
            8'hFF   :  r_t3 = 8'h4F;
        endcase
        end
        
    always@(*)
        begin
        case(w_x[39:32])
            8'h0   :  r_t4 = 8'h70;
            8'h1   :  r_t4 = 8'h2C;
            8'h2   :  r_t4 = 8'hB3;
            8'h3   :  r_t4 = 8'hC0;
            8'h4   :  r_t4 = 8'hE4;
            8'h5   :  r_t4 = 8'h57;
            8'h6   :  r_t4 = 8'hEA;
            8'h7   :  r_t4 = 8'hAE;
            8'h8   :  r_t4 = 8'h23;
            8'h9   :  r_t4 = 8'h6B;
            8'hA   :  r_t4 = 8'h45;
            8'hB   :  r_t4 = 8'hA5;
            8'hC   :  r_t4 = 8'hED;
            8'hD   :  r_t4 = 8'h4F;
            8'hE   :  r_t4 = 8'h1D;
            8'hF   :  r_t4 = 8'h92;
            8'h10   :  r_t4 = 8'h86;
            8'h11   :  r_t4 = 8'hAF;
            8'h12   :  r_t4 = 8'h7C;
            8'h13   :  r_t4 = 8'h1F;
            8'h14   :  r_t4 = 8'h3E;
            8'h15   :  r_t4 = 8'hDC;
            8'h16   :  r_t4 = 8'h5E;
            8'h17   :  r_t4 = 8'hB;
            8'h18   :  r_t4 = 8'hA6;
            8'h19   :  r_t4 = 8'h39;
            8'h1A   :  r_t4 = 8'hD5;
            8'h1B   :  r_t4 = 8'h5D;
            8'h1C   :  r_t4 = 8'hD9;
            8'h1D   :  r_t4 = 8'h5A;
            8'h1E   :  r_t4 = 8'h51;
            8'h1F   :  r_t4 = 8'h6C;
            8'h20   :  r_t4 = 8'h8B;
            8'h21   :  r_t4 = 8'h9A;
            8'h22   :  r_t4 = 8'hFB;
            8'h23   :  r_t4 = 8'hB0;
            8'h24   :  r_t4 = 8'h74;
            8'h25   :  r_t4 = 8'h2B;
            8'h26   :  r_t4 = 8'hF0;
            8'h27   :  r_t4 = 8'h84;
            8'h28   :  r_t4 = 8'hDF;
            8'h29   :  r_t4 = 8'hCB;
            8'h2A   :  r_t4 = 8'h34;
            8'h2B   :  r_t4 = 8'h76;
            8'h2C   :  r_t4 = 8'h6D;
            8'h2D   :  r_t4 = 8'hA9;
            8'h2E   :  r_t4 = 8'hD1;
            8'h2F   :  r_t4 = 8'h4;
            8'h30   :  r_t4 = 8'h14;
            8'h31   :  r_t4 = 8'h3A;
            8'h32   :  r_t4 = 8'hDE;
            8'h33   :  r_t4 = 8'h11;
            8'h34   :  r_t4 = 8'h32;
            8'h35   :  r_t4 = 8'h9C;
            8'h36   :  r_t4 = 8'h53;
            8'h37   :  r_t4 = 8'hF2;
            8'h38   :  r_t4 = 8'hFE;
            8'h39   :  r_t4 = 8'hCF;
            8'h3A   :  r_t4 = 8'hC3;
            8'h3B   :  r_t4 = 8'h7A;
            8'h3C   :  r_t4 = 8'h24;
            8'h3D   :  r_t4 = 8'hE8;
            8'h3E   :  r_t4 = 8'h60;
            8'h3F   :  r_t4 = 8'h69;
            8'h40   :  r_t4 = 8'hAA;
            8'h41   :  r_t4 = 8'hA0;
            8'h42   :  r_t4 = 8'hA1;
            8'h43   :  r_t4 = 8'h62;
            8'h44   :  r_t4 = 8'h54;
            8'h45   :  r_t4 = 8'h1E;
            8'h46   :  r_t4 = 8'hE0;
            8'h47   :  r_t4 = 8'h64;
            8'h48   :  r_t4 = 8'h10;
            8'h49   :  r_t4 = 8'h0;
            8'h4A   :  r_t4 = 8'hA3;
            8'h4B   :  r_t4 = 8'h75;
            8'h4C   :  r_t4 = 8'h8A;
            8'h4D   :  r_t4 = 8'hE6;
            8'h4E   :  r_t4 = 8'h9;
            8'h4F   :  r_t4 = 8'hDD;
            8'h50   :  r_t4 = 8'h87;
            8'h51   :  r_t4 = 8'h83;
            8'h52   :  r_t4 = 8'hCD;
            8'h53   :  r_t4 = 8'h90;
            8'h54   :  r_t4 = 8'h73;
            8'h55   :  r_t4 = 8'hF6;
            8'h56   :  r_t4 = 8'h9D;
            8'h57   :  r_t4 = 8'hBF;
            8'h58   :  r_t4 = 8'h52;
            8'h59   :  r_t4 = 8'hD8;
            8'h5A   :  r_t4 = 8'hC8;
            8'h5B   :  r_t4 = 8'hC6;
            8'h5C   :  r_t4 = 8'h81;
            8'h5D   :  r_t4 = 8'h6F;
            8'h5E   :  r_t4 = 8'h13;
            8'h5F   :  r_t4 = 8'h63;
            8'h60   :  r_t4 = 8'hE9;
            8'h61   :  r_t4 = 8'hA7;
            8'h62   :  r_t4 = 8'h9F;
            8'h63   :  r_t4 = 8'hBC;
            8'h64   :  r_t4 = 8'h29;
            8'h65   :  r_t4 = 8'hF9;
            8'h66   :  r_t4 = 8'h2F;
            8'h67   :  r_t4 = 8'hB4;
            8'h68   :  r_t4 = 8'h78;
            8'h69   :  r_t4 = 8'h6;
            8'h6A   :  r_t4 = 8'hE7;
            8'h6B   :  r_t4 = 8'h71;
            8'h6C   :  r_t4 = 8'hD4;
            8'h6D   :  r_t4 = 8'hAB;
            8'h6E   :  r_t4 = 8'h88;
            8'h6F   :  r_t4 = 8'h8D;
            8'h70   :  r_t4 = 8'h72;
            8'h71   :  r_t4 = 8'hB9;
            8'h72   :  r_t4 = 8'hF8;
            8'h73   :  r_t4 = 8'hAC;
            8'h74   :  r_t4 = 8'h36;
            8'h75   :  r_t4 = 8'h2A;
            8'h76   :  r_t4 = 8'h3C;
            8'h77   :  r_t4 = 8'hF1;
            8'h78   :  r_t4 = 8'h40;
            8'h79   :  r_t4 = 8'hD3;
            8'h7A   :  r_t4 = 8'hBB;
            8'h7B   :  r_t4 = 8'h43;
            8'h7C   :  r_t4 = 8'h15;
            8'h7D   :  r_t4 = 8'hAD;
            8'h7E   :  r_t4 = 8'h77;
            8'h7F   :  r_t4 = 8'h80;
            8'h80   :  r_t4 = 8'h82;
            8'h81   :  r_t4 = 8'hEC;
            8'h82   :  r_t4 = 8'h27;
            8'h83   :  r_t4 = 8'hE5;
            8'h84   :  r_t4 = 8'h85;
            8'h85   :  r_t4 = 8'h35;
            8'h86   :  r_t4 = 8'hC;
            8'h87   :  r_t4 = 8'h41;
            8'h88   :  r_t4 = 8'hEF;
            8'h89   :  r_t4 = 8'h93;
            8'h8A   :  r_t4 = 8'h19;
            8'h8B   :  r_t4 = 8'h21;
            8'h8C   :  r_t4 = 8'hE;
            8'h8D   :  r_t4 = 8'h4E;
            8'h8E   :  r_t4 = 8'h65;
            8'h8F   :  r_t4 = 8'hBD;
            8'h90   :  r_t4 = 8'hB8;
            8'h91   :  r_t4 = 8'h8F;
            8'h92   :  r_t4 = 8'hEB;
            8'h93   :  r_t4 = 8'hCE;
            8'h94   :  r_t4 = 8'h30;
            8'h95   :  r_t4 = 8'h5F;
            8'h96   :  r_t4 = 8'hC5;
            8'h97   :  r_t4 = 8'h1A;
            8'h98   :  r_t4 = 8'hE1;
            8'h99   :  r_t4 = 8'hCA;
            8'h9A   :  r_t4 = 8'h47;
            8'h9B   :  r_t4 = 8'h3D;
            8'h9C   :  r_t4 = 8'h1;
            8'h9D   :  r_t4 = 8'hD6;
            8'h9E   :  r_t4 = 8'h56;
            8'h9F   :  r_t4 = 8'h4D;
            8'hA0   :  r_t4 = 8'hD;
            8'hA1   :  r_t4 = 8'h66;
            8'hA2   :  r_t4 = 8'hCC;
            8'hA3   :  r_t4 = 8'h2D;
            8'hA4   :  r_t4 = 8'h12;
            8'hA5   :  r_t4 = 8'h20;
            8'hA6   :  r_t4 = 8'hB1;
            8'hA7   :  r_t4 = 8'h99;
            8'hA8   :  r_t4 = 8'h4C;
            8'hA9   :  r_t4 = 8'hC2;
            8'hAA   :  r_t4 = 8'h7E;
            8'hAB   :  r_t4 = 8'h5;
            8'hAC   :  r_t4 = 8'hB7;
            8'hAD   :  r_t4 = 8'h31;
            8'hAE   :  r_t4 = 8'h17;
            8'hAF   :  r_t4 = 8'hD7;
            8'hB0   :  r_t4 = 8'h58;
            8'hB1   :  r_t4 = 8'h61;
            8'hB2   :  r_t4 = 8'h1B;
            8'hB3   :  r_t4 = 8'h1C;
            8'hB4   :  r_t4 = 8'hF;
            8'hB5   :  r_t4 = 8'h16;
            8'hB6   :  r_t4 = 8'h18;
            8'hB7   :  r_t4 = 8'h22;
            8'hB8   :  r_t4 = 8'h44;
            8'hB9   :  r_t4 = 8'hB2;
            8'hBA   :  r_t4 = 8'hB5;
            8'hBB   :  r_t4 = 8'h91;
            8'hBC   :  r_t4 = 8'h8;
            8'hBD   :  r_t4 = 8'hA8;
            8'hBE   :  r_t4 = 8'hFC;
            8'hBF   :  r_t4 = 8'h50;
            8'hC0   :  r_t4 = 8'hD0;
            8'hC1   :  r_t4 = 8'h7D;
            8'hC2   :  r_t4 = 8'h89;
            8'hC3   :  r_t4 = 8'h97;
            8'hC4   :  r_t4 = 8'h5B;
            8'hC5   :  r_t4 = 8'h95;
            8'hC6   :  r_t4 = 8'hFF;
            8'hC7   :  r_t4 = 8'hD2;
            8'hC8   :  r_t4 = 8'hC4;
            8'hC9   :  r_t4 = 8'h48;
            8'hCA   :  r_t4 = 8'hF7;
            8'hCB   :  r_t4 = 8'hDB;
            8'hCC   :  r_t4 = 8'h3;
            8'hCD   :  r_t4 = 8'hDA;
            8'hCE   :  r_t4 = 8'h3F;
            8'hCF   :  r_t4 = 8'h94;
            8'hD0   :  r_t4 = 8'h5C;
            8'hD1   :  r_t4 = 8'h2;
            8'hD2   :  r_t4 = 8'h4A;
            8'hD3   :  r_t4 = 8'h33;
            8'hD4   :  r_t4 = 8'h67;
            8'hD5   :  r_t4 = 8'hF3;
            8'hD6   :  r_t4 = 8'h7F;
            8'hD7   :  r_t4 = 8'hE2;
            8'hD8   :  r_t4 = 8'h9B;
            8'hD9   :  r_t4 = 8'h26;
            8'hDA   :  r_t4 = 8'h37;
            8'hDB   :  r_t4 = 8'h3B;
            8'hDC   :  r_t4 = 8'h96;
            8'hDD   :  r_t4 = 8'h4B;
            8'hDE   :  r_t4 = 8'hBE;
            8'hDF   :  r_t4 = 8'h2E;
            8'hE0   :  r_t4 = 8'h79;
            8'hE1   :  r_t4 = 8'h8C;
            8'hE2   :  r_t4 = 8'h6E;
            8'hE3   :  r_t4 = 8'h8E;
            8'hE4   :  r_t4 = 8'hF5;
            8'hE5   :  r_t4 = 8'hB6;
            8'hE6   :  r_t4 = 8'hFD;
            8'hE7   :  r_t4 = 8'h59;
            8'hE8   :  r_t4 = 8'h98;
            8'hE9   :  r_t4 = 8'h6A;
            8'hEA   :  r_t4 = 8'h46;
            8'hEB   :  r_t4 = 8'hBA;
            8'hEC   :  r_t4 = 8'h25;
            8'hED   :  r_t4 = 8'h42;
            8'hEE   :  r_t4 = 8'hA2;
            8'hEF   :  r_t4 = 8'hFA;
            8'hF0   :  r_t4 = 8'h7;
            8'hF1   :  r_t4 = 8'h55;
            8'hF2   :  r_t4 = 8'hEE;
            8'hF3   :  r_t4 = 8'hA;
            8'hF4   :  r_t4 = 8'h49;
            8'hF5   :  r_t4 = 8'h68;
            8'hF6   :  r_t4 = 8'h38;
            8'hF7   :  r_t4 = 8'hA4;
            8'hF8   :  r_t4 = 8'h28;
            8'hF9   :  r_t4 = 8'h7B;
            8'hFA   :  r_t4 = 8'hC9;
            8'hFB   :  r_t4 = 8'hC1;
            8'hFC   :  r_t4 = 8'hE3;
            8'hFD   :  r_t4 = 8'hF4;
            8'hFE   :  r_t4 = 8'hC7;
            8'hFF   :  r_t4 = 8'h9E;
        endcase
        end
        
    always@(*)
        begin
        case(w_x[31:24])
            8'h0   :  r_t5 = 8'hE0;
            8'h1   :  r_t5 = 8'h5;
            8'h2   :  r_t5 = 8'h58;
            8'h3   :  r_t5 = 8'hD9;
            8'h4   :  r_t5 = 8'h67;
            8'h5   :  r_t5 = 8'h4E;
            8'h6   :  r_t5 = 8'h81;
            8'h7   :  r_t5 = 8'hCB;
            8'h8   :  r_t5 = 8'hC9;
            8'h9   :  r_t5 = 8'hB;
            8'hA   :  r_t5 = 8'hAE;
            8'hB   :  r_t5 = 8'h6A;
            8'hC   :  r_t5 = 8'hD5;
            8'hD   :  r_t5 = 8'h18;
            8'hE   :  r_t5 = 8'h5D;
            8'hF   :  r_t5 = 8'h82;
            8'h10   :  r_t5 = 8'h46;
            8'h11   :  r_t5 = 8'hDF;
            8'h12   :  r_t5 = 8'hD6;
            8'h13   :  r_t5 = 8'h27;
            8'h14   :  r_t5 = 8'h8A;
            8'h15   :  r_t5 = 8'h32;
            8'h16   :  r_t5 = 8'h4B;
            8'h17   :  r_t5 = 8'h42;
            8'h18   :  r_t5 = 8'hDB;
            8'h19   :  r_t5 = 8'h1C;
            8'h1A   :  r_t5 = 8'h9E;
            8'h1B   :  r_t5 = 8'h9C;
            8'h1C   :  r_t5 = 8'h3A;
            8'h1D   :  r_t5 = 8'hCA;
            8'h1E   :  r_t5 = 8'h25;
            8'h1F   :  r_t5 = 8'h7B;
            8'h20   :  r_t5 = 8'hD;
            8'h21   :  r_t5 = 8'h71;
            8'h22   :  r_t5 = 8'h5F;
            8'h23   :  r_t5 = 8'h1F;
            8'h24   :  r_t5 = 8'hF8;
            8'h25   :  r_t5 = 8'hD7;
            8'h26   :  r_t5 = 8'h3E;
            8'h27   :  r_t5 = 8'h9D;
            8'h28   :  r_t5 = 8'h7C;
            8'h29   :  r_t5 = 8'h60;
            8'h2A   :  r_t5 = 8'hB9;
            8'h2B   :  r_t5 = 8'hBE;
            8'h2C   :  r_t5 = 8'hBC;
            8'h2D   :  r_t5 = 8'h8B;
            8'h2E   :  r_t5 = 8'h16;
            8'h2F   :  r_t5 = 8'h34;
            8'h30   :  r_t5 = 8'h4D;
            8'h31   :  r_t5 = 8'hC3;
            8'h32   :  r_t5 = 8'h72;
            8'h33   :  r_t5 = 8'h95;
            8'h34   :  r_t5 = 8'hAB;
            8'h35   :  r_t5 = 8'h8E;
            8'h36   :  r_t5 = 8'hBA;
            8'h37   :  r_t5 = 8'h7A;
            8'h38   :  r_t5 = 8'hB3;
            8'h39   :  r_t5 = 8'h2;
            8'h3A   :  r_t5 = 8'hB4;
            8'h3B   :  r_t5 = 8'hAD;
            8'h3C   :  r_t5 = 8'hA2;
            8'h3D   :  r_t5 = 8'hAC;
            8'h3E   :  r_t5 = 8'hD8;
            8'h3F   :  r_t5 = 8'h9A;
            8'h40   :  r_t5 = 8'h17;
            8'h41   :  r_t5 = 8'h1A;
            8'h42   :  r_t5 = 8'h35;
            8'h43   :  r_t5 = 8'hCC;
            8'h44   :  r_t5 = 8'hF7;
            8'h45   :  r_t5 = 8'h99;
            8'h46   :  r_t5 = 8'h61;
            8'h47   :  r_t5 = 8'h5A;
            8'h48   :  r_t5 = 8'hE8;
            8'h49   :  r_t5 = 8'h24;
            8'h4A   :  r_t5 = 8'h56;
            8'h4B   :  r_t5 = 8'h40;
            8'h4C   :  r_t5 = 8'hE1;
            8'h4D   :  r_t5 = 8'h63;
            8'h4E   :  r_t5 = 8'h9;
            8'h4F   :  r_t5 = 8'h33;
            8'h50   :  r_t5 = 8'hBF;
            8'h51   :  r_t5 = 8'h98;
            8'h52   :  r_t5 = 8'h97;
            8'h53   :  r_t5 = 8'h85;
            8'h54   :  r_t5 = 8'h68;
            8'h55   :  r_t5 = 8'hFC;
            8'h56   :  r_t5 = 8'hEC;
            8'h57   :  r_t5 = 8'hA;
            8'h58   :  r_t5 = 8'hDA;
            8'h59   :  r_t5 = 8'h6F;
            8'h5A   :  r_t5 = 8'h53;
            8'h5B   :  r_t5 = 8'h62;
            8'h5C   :  r_t5 = 8'hA3;
            8'h5D   :  r_t5 = 8'h2E;
            8'h5E   :  r_t5 = 8'h8;
            8'h5F   :  r_t5 = 8'hAF;
            8'h60   :  r_t5 = 8'h28;
            8'h61   :  r_t5 = 8'hB0;
            8'h62   :  r_t5 = 8'h74;
            8'h63   :  r_t5 = 8'hC2;
            8'h64   :  r_t5 = 8'hBD;
            8'h65   :  r_t5 = 8'h36;
            8'h66   :  r_t5 = 8'h22;
            8'h67   :  r_t5 = 8'h38;
            8'h68   :  r_t5 = 8'h64;
            8'h69   :  r_t5 = 8'h1E;
            8'h6A   :  r_t5 = 8'h39;
            8'h6B   :  r_t5 = 8'h2C;
            8'h6C   :  r_t5 = 8'hA6;
            8'h6D   :  r_t5 = 8'h30;
            8'h6E   :  r_t5 = 8'hE5;
            8'h6F   :  r_t5 = 8'h44;
            8'h70   :  r_t5 = 8'hFD;
            8'h71   :  r_t5 = 8'h88;
            8'h72   :  r_t5 = 8'h9F;
            8'h73   :  r_t5 = 8'h65;
            8'h74   :  r_t5 = 8'h87;
            8'h75   :  r_t5 = 8'h6B;
            8'h76   :  r_t5 = 8'hF4;
            8'h77   :  r_t5 = 8'h23;
            8'h78   :  r_t5 = 8'h48;
            8'h79   :  r_t5 = 8'h10;
            8'h7A   :  r_t5 = 8'hD1;
            8'h7B   :  r_t5 = 8'h51;
            8'h7C   :  r_t5 = 8'hC0;
            8'h7D   :  r_t5 = 8'hF9;
            8'h7E   :  r_t5 = 8'hD2;
            8'h7F   :  r_t5 = 8'hA0;
            8'h80   :  r_t5 = 8'h55;
            8'h81   :  r_t5 = 8'hA1;
            8'h82   :  r_t5 = 8'h41;
            8'h83   :  r_t5 = 8'hFA;
            8'h84   :  r_t5 = 8'h43;
            8'h85   :  r_t5 = 8'h13;
            8'h86   :  r_t5 = 8'hC4;
            8'h87   :  r_t5 = 8'h2F;
            8'h88   :  r_t5 = 8'hA8;
            8'h89   :  r_t5 = 8'hB6;
            8'h8A   :  r_t5 = 8'h3C;
            8'h8B   :  r_t5 = 8'h2B;
            8'h8C   :  r_t5 = 8'hC1;
            8'h8D   :  r_t5 = 8'hFF;
            8'h8E   :  r_t5 = 8'hC8;
            8'h8F   :  r_t5 = 8'hA5;
            8'h90   :  r_t5 = 8'h20;
            8'h91   :  r_t5 = 8'h89;
            8'h92   :  r_t5 = 8'h0;
            8'h93   :  r_t5 = 8'h90;
            8'h94   :  r_t5 = 8'h47;
            8'h95   :  r_t5 = 8'hEF;
            8'h96   :  r_t5 = 8'hEA;
            8'h97   :  r_t5 = 8'hB7;
            8'h98   :  r_t5 = 8'h15;
            8'h99   :  r_t5 = 8'h6;
            8'h9A   :  r_t5 = 8'hCD;
            8'h9B   :  r_t5 = 8'hB5;
            8'h9C   :  r_t5 = 8'h12;
            8'h9D   :  r_t5 = 8'h7E;
            8'h9E   :  r_t5 = 8'hBB;
            8'h9F   :  r_t5 = 8'h29;
            8'hA0   :  r_t5 = 8'hF;
            8'hA1   :  r_t5 = 8'hB8;
            8'hA2   :  r_t5 = 8'h7;
            8'hA3   :  r_t5 = 8'h4;
            8'hA4   :  r_t5 = 8'h9B;
            8'hA5   :  r_t5 = 8'h94;
            8'hA6   :  r_t5 = 8'h21;
            8'hA7   :  r_t5 = 8'h66;
            8'hA8   :  r_t5 = 8'hE6;
            8'hA9   :  r_t5 = 8'hCE;
            8'hAA   :  r_t5 = 8'hED;
            8'hAB   :  r_t5 = 8'hE7;
            8'hAC   :  r_t5 = 8'h3B;
            8'hAD   :  r_t5 = 8'hFE;
            8'hAE   :  r_t5 = 8'h7F;
            8'hAF   :  r_t5 = 8'hC5;
            8'hB0   :  r_t5 = 8'hA4;
            8'hB1   :  r_t5 = 8'h37;
            8'hB2   :  r_t5 = 8'hB1;
            8'hB3   :  r_t5 = 8'h4C;
            8'hB4   :  r_t5 = 8'h91;
            8'hB5   :  r_t5 = 8'h6E;
            8'hB6   :  r_t5 = 8'h8D;
            8'hB7   :  r_t5 = 8'h76;
            8'hB8   :  r_t5 = 8'h3;
            8'hB9   :  r_t5 = 8'h2D;
            8'hBA   :  r_t5 = 8'hDE;
            8'hBB   :  r_t5 = 8'h96;
            8'hBC   :  r_t5 = 8'h26;
            8'hBD   :  r_t5 = 8'h7D;
            8'hBE   :  r_t5 = 8'hC6;
            8'hBF   :  r_t5 = 8'h5C;
            8'hC0   :  r_t5 = 8'hD3;
            8'hC1   :  r_t5 = 8'hF2;
            8'hC2   :  r_t5 = 8'h4F;
            8'hC3   :  r_t5 = 8'h19;
            8'hC4   :  r_t5 = 8'h3F;
            8'hC5   :  r_t5 = 8'hDC;
            8'hC6   :  r_t5 = 8'h79;
            8'hC7   :  r_t5 = 8'h1D;
            8'hC8   :  r_t5 = 8'h52;
            8'hC9   :  r_t5 = 8'hEB;
            8'hCA   :  r_t5 = 8'hF3;
            8'hCB   :  r_t5 = 8'h6D;
            8'hCC   :  r_t5 = 8'h5E;
            8'hCD   :  r_t5 = 8'hFB;
            8'hCE   :  r_t5 = 8'h69;
            8'hCF   :  r_t5 = 8'hB2;
            8'hD0   :  r_t5 = 8'hF0;
            8'hD1   :  r_t5 = 8'h31;
            8'hD2   :  r_t5 = 8'hC;
            8'hD3   :  r_t5 = 8'hD4;
            8'hD4   :  r_t5 = 8'hCF;
            8'hD5   :  r_t5 = 8'h8C;
            8'hD6   :  r_t5 = 8'hE2;
            8'hD7   :  r_t5 = 8'h75;
            8'hD8   :  r_t5 = 8'hA9;
            8'hD9   :  r_t5 = 8'h4A;
            8'hDA   :  r_t5 = 8'h57;
            8'hDB   :  r_t5 = 8'h84;
            8'hDC   :  r_t5 = 8'h11;
            8'hDD   :  r_t5 = 8'h45;
            8'hDE   :  r_t5 = 8'h1B;
            8'hDF   :  r_t5 = 8'hF5;
            8'hE0   :  r_t5 = 8'hE4;
            8'hE1   :  r_t5 = 8'hE;
            8'hE2   :  r_t5 = 8'h73;
            8'hE3   :  r_t5 = 8'hAA;
            8'hE4   :  r_t5 = 8'hF1;
            8'hE5   :  r_t5 = 8'hDD;
            8'hE6   :  r_t5 = 8'h59;
            8'hE7   :  r_t5 = 8'h14;
            8'hE8   :  r_t5 = 8'h6C;
            8'hE9   :  r_t5 = 8'h92;
            8'hEA   :  r_t5 = 8'h54;
            8'hEB   :  r_t5 = 8'hD0;
            8'hEC   :  r_t5 = 8'h78;
            8'hED   :  r_t5 = 8'h70;
            8'hEE   :  r_t5 = 8'hE3;
            8'hEF   :  r_t5 = 8'h49;
            8'hF0   :  r_t5 = 8'h80;
            8'hF1   :  r_t5 = 8'h50;
            8'hF2   :  r_t5 = 8'hA7;
            8'hF3   :  r_t5 = 8'hF6;
            8'hF4   :  r_t5 = 8'h77;
            8'hF5   :  r_t5 = 8'h93;
            8'hF6   :  r_t5 = 8'h86;
            8'hF7   :  r_t5 = 8'h83;
            8'hF8   :  r_t5 = 8'h2A;
            8'hF9   :  r_t5 = 8'hC7;
            8'hFA   :  r_t5 = 8'h5B;
            8'hFB   :  r_t5 = 8'hE9;
            8'hFC   :  r_t5 = 8'hEE;
            8'hFD   :  r_t5 = 8'h8F;
            8'hFE   :  r_t5 = 8'h1;
            8'hFF   :  r_t5 = 8'h3D;
        endcase
        end
        
    always@(*)
        begin
        case(w_x[23:16])
            8'h0   :  r_t6 = 8'h38;
            8'h1   :  r_t6 = 8'h41;
            8'h2   :  r_t6 = 8'h16;
            8'h3   :  r_t6 = 8'h76;
            8'h4   :  r_t6 = 8'hD9;
            8'h5   :  r_t6 = 8'h93;
            8'h6   :  r_t6 = 8'h60;
            8'h7   :  r_t6 = 8'hF2;
            8'h8   :  r_t6 = 8'h72;
            8'h9   :  r_t6 = 8'hC2;
            8'hA   :  r_t6 = 8'hAB;
            8'hB   :  r_t6 = 8'h9A;
            8'hC   :  r_t6 = 8'h75;
            8'hD   :  r_t6 = 8'h6;
            8'hE   :  r_t6 = 8'h57;
            8'hF   :  r_t6 = 8'hA0;
            8'h10   :  r_t6 = 8'h91;
            8'h11   :  r_t6 = 8'hF7;
            8'h12   :  r_t6 = 8'hB5;
            8'h13   :  r_t6 = 8'hC9;
            8'h14   :  r_t6 = 8'hA2;
            8'h15   :  r_t6 = 8'h8C;
            8'h16   :  r_t6 = 8'hD2;
            8'h17   :  r_t6 = 8'h90;
            8'h18   :  r_t6 = 8'hF6;
            8'h19   :  r_t6 = 8'h7;
            8'h1A   :  r_t6 = 8'hA7;
            8'h1B   :  r_t6 = 8'h27;
            8'h1C   :  r_t6 = 8'h8E;
            8'h1D   :  r_t6 = 8'hB2;
            8'h1E   :  r_t6 = 8'h49;
            8'h1F   :  r_t6 = 8'hDE;
            8'h20   :  r_t6 = 8'h43;
            8'h21   :  r_t6 = 8'h5C;
            8'h22   :  r_t6 = 8'hD7;
            8'h23   :  r_t6 = 8'hC7;
            8'h24   :  r_t6 = 8'h3E;
            8'h25   :  r_t6 = 8'hF5;
            8'h26   :  r_t6 = 8'h8F;
            8'h27   :  r_t6 = 8'h67;
            8'h28   :  r_t6 = 8'h1F;
            8'h29   :  r_t6 = 8'h18;
            8'h2A   :  r_t6 = 8'h6E;
            8'h2B   :  r_t6 = 8'hAF;
            8'h2C   :  r_t6 = 8'h2F;
            8'h2D   :  r_t6 = 8'hE2;
            8'h2E   :  r_t6 = 8'h85;
            8'h2F   :  r_t6 = 8'hD;
            8'h30   :  r_t6 = 8'h53;
            8'h31   :  r_t6 = 8'hF0;
            8'h32   :  r_t6 = 8'h9C;
            8'h33   :  r_t6 = 8'h65;
            8'h34   :  r_t6 = 8'hEA;
            8'h35   :  r_t6 = 8'hA3;
            8'h36   :  r_t6 = 8'hAE;
            8'h37   :  r_t6 = 8'h9E;
            8'h38   :  r_t6 = 8'hEC;
            8'h39   :  r_t6 = 8'h80;
            8'h3A   :  r_t6 = 8'h2D;
            8'h3B   :  r_t6 = 8'h6B;
            8'h3C   :  r_t6 = 8'hA8;
            8'h3D   :  r_t6 = 8'h2B;
            8'h3E   :  r_t6 = 8'h36;
            8'h3F   :  r_t6 = 8'hA6;
            8'h40   :  r_t6 = 8'hC5;
            8'h41   :  r_t6 = 8'h86;
            8'h42   :  r_t6 = 8'h4D;
            8'h43   :  r_t6 = 8'h33;
            8'h44   :  r_t6 = 8'hFD;
            8'h45   :  r_t6 = 8'h66;
            8'h46   :  r_t6 = 8'h58;
            8'h47   :  r_t6 = 8'h96;
            8'h48   :  r_t6 = 8'h3A;
            8'h49   :  r_t6 = 8'h9;
            8'h4A   :  r_t6 = 8'h95;
            8'h4B   :  r_t6 = 8'h10;
            8'h4C   :  r_t6 = 8'h78;
            8'h4D   :  r_t6 = 8'hD8;
            8'h4E   :  r_t6 = 8'h42;
            8'h4F   :  r_t6 = 8'hCC;
            8'h50   :  r_t6 = 8'hEF;
            8'h51   :  r_t6 = 8'h26;
            8'h52   :  r_t6 = 8'hE5;
            8'h53   :  r_t6 = 8'h61;
            8'h54   :  r_t6 = 8'h1A;
            8'h55   :  r_t6 = 8'h3F;
            8'h56   :  r_t6 = 8'h3B;
            8'h57   :  r_t6 = 8'h82;
            8'h58   :  r_t6 = 8'hB6;
            8'h59   :  r_t6 = 8'hDB;
            8'h5A   :  r_t6 = 8'hD4;
            8'h5B   :  r_t6 = 8'h98;
            8'h5C   :  r_t6 = 8'hE8;
            8'h5D   :  r_t6 = 8'h8B;
            8'h5E   :  r_t6 = 8'h2;
            8'h5F   :  r_t6 = 8'hEB;
            8'h60   :  r_t6 = 8'hA;
            8'h61   :  r_t6 = 8'h2C;
            8'h62   :  r_t6 = 8'h1D;
            8'h63   :  r_t6 = 8'hB0;
            8'h64   :  r_t6 = 8'h6F;
            8'h65   :  r_t6 = 8'h8D;
            8'h66   :  r_t6 = 8'h88;
            8'h67   :  r_t6 = 8'hE;
            8'h68   :  r_t6 = 8'h19;
            8'h69   :  r_t6 = 8'h87;
            8'h6A   :  r_t6 = 8'h4E;
            8'h6B   :  r_t6 = 8'hB;
            8'h6C   :  r_t6 = 8'hA9;
            8'h6D   :  r_t6 = 8'hC;
            8'h6E   :  r_t6 = 8'h79;
            8'h6F   :  r_t6 = 8'h11;
            8'h70   :  r_t6 = 8'h7F;
            8'h71   :  r_t6 = 8'h22;
            8'h72   :  r_t6 = 8'hE7;
            8'h73   :  r_t6 = 8'h59;
            8'h74   :  r_t6 = 8'hE1;
            8'h75   :  r_t6 = 8'hDA;
            8'h76   :  r_t6 = 8'h3D;
            8'h77   :  r_t6 = 8'hC8;
            8'h78   :  r_t6 = 8'h12;
            8'h79   :  r_t6 = 8'h4;
            8'h7A   :  r_t6 = 8'h74;
            8'h7B   :  r_t6 = 8'h54;
            8'h7C   :  r_t6 = 8'h30;
            8'h7D   :  r_t6 = 8'h7E;
            8'h7E   :  r_t6 = 8'hB4;
            8'h7F   :  r_t6 = 8'h28;
            8'h80   :  r_t6 = 8'h55;
            8'h81   :  r_t6 = 8'h68;
            8'h82   :  r_t6 = 8'h50;
            8'h83   :  r_t6 = 8'hBE;
            8'h84   :  r_t6 = 8'hD0;
            8'h85   :  r_t6 = 8'hC4;
            8'h86   :  r_t6 = 8'h31;
            8'h87   :  r_t6 = 8'hCB;
            8'h88   :  r_t6 = 8'h2A;
            8'h89   :  r_t6 = 8'hAD;
            8'h8A   :  r_t6 = 8'hF;
            8'h8B   :  r_t6 = 8'hCA;
            8'h8C   :  r_t6 = 8'h70;
            8'h8D   :  r_t6 = 8'hFF;
            8'h8E   :  r_t6 = 8'h32;
            8'h8F   :  r_t6 = 8'h69;
            8'h90   :  r_t6 = 8'h8;
            8'h91   :  r_t6 = 8'h62;
            8'h92   :  r_t6 = 8'h0;
            8'h93   :  r_t6 = 8'h24;
            8'h94   :  r_t6 = 8'hD1;
            8'h95   :  r_t6 = 8'hFB;
            8'h96   :  r_t6 = 8'hBA;
            8'h97   :  r_t6 = 8'hED;
            8'h98   :  r_t6 = 8'h45;
            8'h99   :  r_t6 = 8'h81;
            8'h9A   :  r_t6 = 8'h73;
            8'h9B   :  r_t6 = 8'h6D;
            8'h9C   :  r_t6 = 8'h84;
            8'h9D   :  r_t6 = 8'h9F;
            8'h9E   :  r_t6 = 8'hEE;
            8'h9F   :  r_t6 = 8'h4A;
            8'hA0   :  r_t6 = 8'hC3;
            8'hA1   :  r_t6 = 8'h2E;
            8'hA2   :  r_t6 = 8'hC1;
            8'hA3   :  r_t6 = 8'h1;
            8'hA4   :  r_t6 = 8'hE6;
            8'hA5   :  r_t6 = 8'h25;
            8'hA6   :  r_t6 = 8'h48;
            8'hA7   :  r_t6 = 8'h99;
            8'hA8   :  r_t6 = 8'hB9;
            8'hA9   :  r_t6 = 8'hB3;
            8'hAA   :  r_t6 = 8'h7B;
            8'hAB   :  r_t6 = 8'hF9;
            8'hAC   :  r_t6 = 8'hCE;
            8'hAD   :  r_t6 = 8'hBF;
            8'hAE   :  r_t6 = 8'hDF;
            8'hAF   :  r_t6 = 8'h71;
            8'hB0   :  r_t6 = 8'h29;
            8'hB1   :  r_t6 = 8'hCD;
            8'hB2   :  r_t6 = 8'h6C;
            8'hB3   :  r_t6 = 8'h13;
            8'hB4   :  r_t6 = 8'h64;
            8'hB5   :  r_t6 = 8'h9B;
            8'hB6   :  r_t6 = 8'h63;
            8'hB7   :  r_t6 = 8'h9D;
            8'hB8   :  r_t6 = 8'hC0;
            8'hB9   :  r_t6 = 8'h4B;
            8'hBA   :  r_t6 = 8'hB7;
            8'hBB   :  r_t6 = 8'hA5;
            8'hBC   :  r_t6 = 8'h89;
            8'hBD   :  r_t6 = 8'h5F;
            8'hBE   :  r_t6 = 8'hB1;
            8'hBF   :  r_t6 = 8'h17;
            8'hC0   :  r_t6 = 8'hF4;
            8'hC1   :  r_t6 = 8'hBC;
            8'hC2   :  r_t6 = 8'hD3;
            8'hC3   :  r_t6 = 8'h46;
            8'hC4   :  r_t6 = 8'hCF;
            8'hC5   :  r_t6 = 8'h37;
            8'hC6   :  r_t6 = 8'h5E;
            8'hC7   :  r_t6 = 8'h47;
            8'hC8   :  r_t6 = 8'h94;
            8'hC9   :  r_t6 = 8'hFA;
            8'hCA   :  r_t6 = 8'hFC;
            8'hCB   :  r_t6 = 8'h5B;
            8'hCC   :  r_t6 = 8'h97;
            8'hCD   :  r_t6 = 8'hFE;
            8'hCE   :  r_t6 = 8'h5A;
            8'hCF   :  r_t6 = 8'hAC;
            8'hD0   :  r_t6 = 8'h3C;
            8'hD1   :  r_t6 = 8'h4C;
            8'hD2   :  r_t6 = 8'h3;
            8'hD3   :  r_t6 = 8'h35;
            8'hD4   :  r_t6 = 8'hF3;
            8'hD5   :  r_t6 = 8'h23;
            8'hD6   :  r_t6 = 8'hB8;
            8'hD7   :  r_t6 = 8'h5D;
            8'hD8   :  r_t6 = 8'h6A;
            8'hD9   :  r_t6 = 8'h92;
            8'hDA   :  r_t6 = 8'hD5;
            8'hDB   :  r_t6 = 8'h21;
            8'hDC   :  r_t6 = 8'h44;
            8'hDD   :  r_t6 = 8'h51;
            8'hDE   :  r_t6 = 8'hC6;
            8'hDF   :  r_t6 = 8'h7D;
            8'hE0   :  r_t6 = 8'h39;
            8'hE1   :  r_t6 = 8'h83;
            8'hE2   :  r_t6 = 8'hDC;
            8'hE3   :  r_t6 = 8'hAA;
            8'hE4   :  r_t6 = 8'h7C;
            8'hE5   :  r_t6 = 8'h77;
            8'hE6   :  r_t6 = 8'h56;
            8'hE7   :  r_t6 = 8'h5;
            8'hE8   :  r_t6 = 8'h1B;
            8'hE9   :  r_t6 = 8'hA4;
            8'hEA   :  r_t6 = 8'h15;
            8'hEB   :  r_t6 = 8'h34;
            8'hEC   :  r_t6 = 8'h1E;
            8'hED   :  r_t6 = 8'h1C;
            8'hEE   :  r_t6 = 8'hF8;
            8'hEF   :  r_t6 = 8'h52;
            8'hF0   :  r_t6 = 8'h20;
            8'hF1   :  r_t6 = 8'h14;
            8'hF2   :  r_t6 = 8'hE9;
            8'hF3   :  r_t6 = 8'hBD;
            8'hF4   :  r_t6 = 8'hDD;
            8'hF5   :  r_t6 = 8'hE4;
            8'hF6   :  r_t6 = 8'hA1;
            8'hF7   :  r_t6 = 8'hE0;
            8'hF8   :  r_t6 = 8'h8A;
            8'hF9   :  r_t6 = 8'hF1;
            8'hFA   :  r_t6 = 8'hD6;
            8'hFB   :  r_t6 = 8'h7A;
            8'hFC   :  r_t6 = 8'hBB;
            8'hFD   :  r_t6 = 8'hE3;
            8'hFE   :  r_t6 = 8'h40;
            8'hFF   :  r_t6 = 8'h4F;
        endcase
        end
        
    always@(*)
        begin
        case(w_x[15:8])
            8'h0   :  r_t7 = 8'h70;
            8'h1   :  r_t7 = 8'h2C;
            8'h2   :  r_t7 = 8'hB3;
            8'h3   :  r_t7 = 8'hC0;
            8'h4   :  r_t7 = 8'hE4;
            8'h5   :  r_t7 = 8'h57;
            8'h6   :  r_t7 = 8'hEA;
            8'h7   :  r_t7 = 8'hAE;
            8'h8   :  r_t7 = 8'h23;
            8'h9   :  r_t7 = 8'h6B;
            8'hA   :  r_t7 = 8'h45;
            8'hB   :  r_t7 = 8'hA5;
            8'hC   :  r_t7 = 8'hED;
            8'hD   :  r_t7 = 8'h4F;
            8'hE   :  r_t7 = 8'h1D;
            8'hF   :  r_t7 = 8'h92;
            8'h10   :  r_t7 = 8'h86;
            8'h11   :  r_t7 = 8'hAF;
            8'h12   :  r_t7 = 8'h7C;
            8'h13   :  r_t7 = 8'h1F;
            8'h14   :  r_t7 = 8'h3E;
            8'h15   :  r_t7 = 8'hDC;
            8'h16   :  r_t7 = 8'h5E;
            8'h17   :  r_t7 = 8'hB;
            8'h18   :  r_t7 = 8'hA6;
            8'h19   :  r_t7 = 8'h39;
            8'h1A   :  r_t7 = 8'hD5;
            8'h1B   :  r_t7 = 8'h5D;
            8'h1C   :  r_t7 = 8'hD9;
            8'h1D   :  r_t7 = 8'h5A;
            8'h1E   :  r_t7 = 8'h51;
            8'h1F   :  r_t7 = 8'h6C;
            8'h20   :  r_t7 = 8'h8B;
            8'h21   :  r_t7 = 8'h9A;
            8'h22   :  r_t7 = 8'hFB;
            8'h23   :  r_t7 = 8'hB0;
            8'h24   :  r_t7 = 8'h74;
            8'h25   :  r_t7 = 8'h2B;
            8'h26   :  r_t7 = 8'hF0;
            8'h27   :  r_t7 = 8'h84;
            8'h28   :  r_t7 = 8'hDF;
            8'h29   :  r_t7 = 8'hCB;
            8'h2A   :  r_t7 = 8'h34;
            8'h2B   :  r_t7 = 8'h76;
            8'h2C   :  r_t7 = 8'h6D;
            8'h2D   :  r_t7 = 8'hA9;
            8'h2E   :  r_t7 = 8'hD1;
            8'h2F   :  r_t7 = 8'h4;
            8'h30   :  r_t7 = 8'h14;
            8'h31   :  r_t7 = 8'h3A;
            8'h32   :  r_t7 = 8'hDE;
            8'h33   :  r_t7 = 8'h11;
            8'h34   :  r_t7 = 8'h32;
            8'h35   :  r_t7 = 8'h9C;
            8'h36   :  r_t7 = 8'h53;
            8'h37   :  r_t7 = 8'hF2;
            8'h38   :  r_t7 = 8'hFE;
            8'h39   :  r_t7 = 8'hCF;
            8'h3A   :  r_t7 = 8'hC3;
            8'h3B   :  r_t7 = 8'h7A;
            8'h3C   :  r_t7 = 8'h24;
            8'h3D   :  r_t7 = 8'hE8;
            8'h3E   :  r_t7 = 8'h60;
            8'h3F   :  r_t7 = 8'h69;
            8'h40   :  r_t7 = 8'hAA;
            8'h41   :  r_t7 = 8'hA0;
            8'h42   :  r_t7 = 8'hA1;
            8'h43   :  r_t7 = 8'h62;
            8'h44   :  r_t7 = 8'h54;
            8'h45   :  r_t7 = 8'h1E;
            8'h46   :  r_t7 = 8'hE0;
            8'h47   :  r_t7 = 8'h64;
            8'h48   :  r_t7 = 8'h10;
            8'h49   :  r_t7 = 8'h0;
            8'h4A   :  r_t7 = 8'hA3;
            8'h4B   :  r_t7 = 8'h75;
            8'h4C   :  r_t7 = 8'h8A;
            8'h4D   :  r_t7 = 8'hE6;
            8'h4E   :  r_t7 = 8'h9;
            8'h4F   :  r_t7 = 8'hDD;
            8'h50   :  r_t7 = 8'h87;
            8'h51   :  r_t7 = 8'h83;
            8'h52   :  r_t7 = 8'hCD;
            8'h53   :  r_t7 = 8'h90;
            8'h54   :  r_t7 = 8'h73;
            8'h55   :  r_t7 = 8'hF6;
            8'h56   :  r_t7 = 8'h9D;
            8'h57   :  r_t7 = 8'hBF;
            8'h58   :  r_t7 = 8'h52;
            8'h59   :  r_t7 = 8'hD8;
            8'h5A   :  r_t7 = 8'hC8;
            8'h5B   :  r_t7 = 8'hC6;
            8'h5C   :  r_t7 = 8'h81;
            8'h5D   :  r_t7 = 8'h6F;
            8'h5E   :  r_t7 = 8'h13;
            8'h5F   :  r_t7 = 8'h63;
            8'h60   :  r_t7 = 8'hE9;
            8'h61   :  r_t7 = 8'hA7;
            8'h62   :  r_t7 = 8'h9F;
            8'h63   :  r_t7 = 8'hBC;
            8'h64   :  r_t7 = 8'h29;
            8'h65   :  r_t7 = 8'hF9;
            8'h66   :  r_t7 = 8'h2F;
            8'h67   :  r_t7 = 8'hB4;
            8'h68   :  r_t7 = 8'h78;
            8'h69   :  r_t7 = 8'h6;
            8'h6A   :  r_t7 = 8'hE7;
            8'h6B   :  r_t7 = 8'h71;
            8'h6C   :  r_t7 = 8'hD4;
            8'h6D   :  r_t7 = 8'hAB;
            8'h6E   :  r_t7 = 8'h88;
            8'h6F   :  r_t7 = 8'h8D;
            8'h70   :  r_t7 = 8'h72;
            8'h71   :  r_t7 = 8'hB9;
            8'h72   :  r_t7 = 8'hF8;
            8'h73   :  r_t7 = 8'hAC;
            8'h74   :  r_t7 = 8'h36;
            8'h75   :  r_t7 = 8'h2A;
            8'h76   :  r_t7 = 8'h3C;
            8'h77   :  r_t7 = 8'hF1;
            8'h78   :  r_t7 = 8'h40;
            8'h79   :  r_t7 = 8'hD3;
            8'h7A   :  r_t7 = 8'hBB;
            8'h7B   :  r_t7 = 8'h43;
            8'h7C   :  r_t7 = 8'h15;
            8'h7D   :  r_t7 = 8'hAD;
            8'h7E   :  r_t7 = 8'h77;
            8'h7F   :  r_t7 = 8'h80;
            8'h80   :  r_t7 = 8'h82;
            8'h81   :  r_t7 = 8'hEC;
            8'h82   :  r_t7 = 8'h27;
            8'h83   :  r_t7 = 8'hE5;
            8'h84   :  r_t7 = 8'h85;
            8'h85   :  r_t7 = 8'h35;
            8'h86   :  r_t7 = 8'hC;
            8'h87   :  r_t7 = 8'h41;
            8'h88   :  r_t7 = 8'hEF;
            8'h89   :  r_t7 = 8'h93;
            8'h8A   :  r_t7 = 8'h19;
            8'h8B   :  r_t7 = 8'h21;
            8'h8C   :  r_t7 = 8'hE;
            8'h8D   :  r_t7 = 8'h4E;
            8'h8E   :  r_t7 = 8'h65;
            8'h8F   :  r_t7 = 8'hBD;
            8'h90   :  r_t7 = 8'hB8;
            8'h91   :  r_t7 = 8'h8F;
            8'h92   :  r_t7 = 8'hEB;
            8'h93   :  r_t7 = 8'hCE;
            8'h94   :  r_t7 = 8'h30;
            8'h95   :  r_t7 = 8'h5F;
            8'h96   :  r_t7 = 8'hC5;
            8'h97   :  r_t7 = 8'h1A;
            8'h98   :  r_t7 = 8'hE1;
            8'h99   :  r_t7 = 8'hCA;
            8'h9A   :  r_t7 = 8'h47;
            8'h9B   :  r_t7 = 8'h3D;
            8'h9C   :  r_t7 = 8'h1;
            8'h9D   :  r_t7 = 8'hD6;
            8'h9E   :  r_t7 = 8'h56;
            8'h9F   :  r_t7 = 8'h4D;
            8'hA0   :  r_t7 = 8'hD;
            8'hA1   :  r_t7 = 8'h66;
            8'hA2   :  r_t7 = 8'hCC;
            8'hA3   :  r_t7 = 8'h2D;
            8'hA4   :  r_t7 = 8'h12;
            8'hA5   :  r_t7 = 8'h20;
            8'hA6   :  r_t7 = 8'hB1;
            8'hA7   :  r_t7 = 8'h99;
            8'hA8   :  r_t7 = 8'h4C;
            8'hA9   :  r_t7 = 8'hC2;
            8'hAA   :  r_t7 = 8'h7E;
            8'hAB   :  r_t7 = 8'h5;
            8'hAC   :  r_t7 = 8'hB7;
            8'hAD   :  r_t7 = 8'h31;
            8'hAE   :  r_t7 = 8'h17;
            8'hAF   :  r_t7 = 8'hD7;
            8'hB0   :  r_t7 = 8'h58;
            8'hB1   :  r_t7 = 8'h61;
            8'hB2   :  r_t7 = 8'h1B;
            8'hB3   :  r_t7 = 8'h1C;
            8'hB4   :  r_t7 = 8'hF;
            8'hB5   :  r_t7 = 8'h16;
            8'hB6   :  r_t7 = 8'h18;
            8'hB7   :  r_t7 = 8'h22;
            8'hB8   :  r_t7 = 8'h44;
            8'hB9   :  r_t7 = 8'hB2;
            8'hBA   :  r_t7 = 8'hB5;
            8'hBB   :  r_t7 = 8'h91;
            8'hBC   :  r_t7 = 8'h8;
            8'hBD   :  r_t7 = 8'hA8;
            8'hBE   :  r_t7 = 8'hFC;
            8'hBF   :  r_t7 = 8'h50;
            8'hC0   :  r_t7 = 8'hD0;
            8'hC1   :  r_t7 = 8'h7D;
            8'hC2   :  r_t7 = 8'h89;
            8'hC3   :  r_t7 = 8'h97;
            8'hC4   :  r_t7 = 8'h5B;
            8'hC5   :  r_t7 = 8'h95;
            8'hC6   :  r_t7 = 8'hFF;
            8'hC7   :  r_t7 = 8'hD2;
            8'hC8   :  r_t7 = 8'hC4;
            8'hC9   :  r_t7 = 8'h48;
            8'hCA   :  r_t7 = 8'hF7;
            8'hCB   :  r_t7 = 8'hDB;
            8'hCC   :  r_t7 = 8'h3;
            8'hCD   :  r_t7 = 8'hDA;
            8'hCE   :  r_t7 = 8'h3F;
            8'hCF   :  r_t7 = 8'h94;
            8'hD0   :  r_t7 = 8'h5C;
            8'hD1   :  r_t7 = 8'h2;
            8'hD2   :  r_t7 = 8'h4A;
            8'hD3   :  r_t7 = 8'h33;
            8'hD4   :  r_t7 = 8'h67;
            8'hD5   :  r_t7 = 8'hF3;
            8'hD6   :  r_t7 = 8'h7F;
            8'hD7   :  r_t7 = 8'hE2;
            8'hD8   :  r_t7 = 8'h9B;
            8'hD9   :  r_t7 = 8'h26;
            8'hDA   :  r_t7 = 8'h37;
            8'hDB   :  r_t7 = 8'h3B;
            8'hDC   :  r_t7 = 8'h96;
            8'hDD   :  r_t7 = 8'h4B;
            8'hDE   :  r_t7 = 8'hBE;
            8'hDF   :  r_t7 = 8'h2E;
            8'hE0   :  r_t7 = 8'h79;
            8'hE1   :  r_t7 = 8'h8C;
            8'hE2   :  r_t7 = 8'h6E;
            8'hE3   :  r_t7 = 8'h8E;
            8'hE4   :  r_t7 = 8'hF5;
            8'hE5   :  r_t7 = 8'hB6;
            8'hE6   :  r_t7 = 8'hFD;
            8'hE7   :  r_t7 = 8'h59;
            8'hE8   :  r_t7 = 8'h98;
            8'hE9   :  r_t7 = 8'h6A;
            8'hEA   :  r_t7 = 8'h46;
            8'hEB   :  r_t7 = 8'hBA;
            8'hEC   :  r_t7 = 8'h25;
            8'hED   :  r_t7 = 8'h42;
            8'hEE   :  r_t7 = 8'hA2;
            8'hEF   :  r_t7 = 8'hFA;
            8'hF0   :  r_t7 = 8'h7;
            8'hF1   :  r_t7 = 8'h55;
            8'hF2   :  r_t7 = 8'hEE;
            8'hF3   :  r_t7 = 8'hA;
            8'hF4   :  r_t7 = 8'h49;
            8'hF5   :  r_t7 = 8'h68;
            8'hF6   :  r_t7 = 8'h38;
            8'hF7   :  r_t7 = 8'hA4;
            8'hF8   :  r_t7 = 8'h28;
            8'hF9   :  r_t7 = 8'h7B;
            8'hFA   :  r_t7 = 8'hC9;
            8'hFB   :  r_t7 = 8'hC1;
            8'hFC   :  r_t7 = 8'hE3;
            8'hFD   :  r_t7 = 8'hF4;
            8'hFE   :  r_t7 = 8'hC7;
            8'hFF   :  r_t7 = 8'h9E;
        endcase
        end
        
    always@(*)
        begin
        case(w_x[7:0])
            8'h0   :  r_t8 = 8'h70;
            8'h1   :  r_t8 = 8'h82;
            8'h2   :  r_t8 = 8'h2C;
            8'h3   :  r_t8 = 8'hEC;
            8'h4   :  r_t8 = 8'hB3;
            8'h5   :  r_t8 = 8'h27;
            8'h6   :  r_t8 = 8'hC0;
            8'h7   :  r_t8 = 8'hE5;
            8'h8   :  r_t8 = 8'hE4;
            8'h9   :  r_t8 = 8'h85;
            8'hA   :  r_t8 = 8'h57;
            8'hB   :  r_t8 = 8'h35;
            8'hC   :  r_t8 = 8'hEA;
            8'hD   :  r_t8 = 8'hC;
            8'hE   :  r_t8 = 8'hAE;
            8'hF   :  r_t8 = 8'h41;
            8'h10   :  r_t8 = 8'h23;
            8'h11   :  r_t8 = 8'hEF;
            8'h12   :  r_t8 = 8'h6B;
            8'h13   :  r_t8 = 8'h93;
            8'h14   :  r_t8 = 8'h45;
            8'h15   :  r_t8 = 8'h19;
            8'h16   :  r_t8 = 8'hA5;
            8'h17   :  r_t8 = 8'h21;
            8'h18   :  r_t8 = 8'hED;
            8'h19   :  r_t8 = 8'hE;
            8'h1A   :  r_t8 = 8'h4F;
            8'h1B   :  r_t8 = 8'h4E;
            8'h1C   :  r_t8 = 8'h1D;
            8'h1D   :  r_t8 = 8'h65;
            8'h1E   :  r_t8 = 8'h92;
            8'h1F   :  r_t8 = 8'hBD;
            8'h20   :  r_t8 = 8'h86;
            8'h21   :  r_t8 = 8'hB8;
            8'h22   :  r_t8 = 8'hAF;
            8'h23   :  r_t8 = 8'h8F;
            8'h24   :  r_t8 = 8'h7C;
            8'h25   :  r_t8 = 8'hEB;
            8'h26   :  r_t8 = 8'h1F;
            8'h27   :  r_t8 = 8'hCE;
            8'h28   :  r_t8 = 8'h3E;
            8'h29   :  r_t8 = 8'h30;
            8'h2A   :  r_t8 = 8'hDC;
            8'h2B   :  r_t8 = 8'h5F;
            8'h2C   :  r_t8 = 8'h5E;
            8'h2D   :  r_t8 = 8'hC5;
            8'h2E   :  r_t8 = 8'hB;
            8'h2F   :  r_t8 = 8'h1A;
            8'h30   :  r_t8 = 8'hA6;
            8'h31   :  r_t8 = 8'hE1;
            8'h32   :  r_t8 = 8'h39;
            8'h33   :  r_t8 = 8'hCA;
            8'h34   :  r_t8 = 8'hD5;
            8'h35   :  r_t8 = 8'h47;
            8'h36   :  r_t8 = 8'h5D;
            8'h37   :  r_t8 = 8'h3D;
            8'h38   :  r_t8 = 8'hD9;
            8'h39   :  r_t8 = 8'h1;
            8'h3A   :  r_t8 = 8'h5A;
            8'h3B   :  r_t8 = 8'hD6;
            8'h3C   :  r_t8 = 8'h51;
            8'h3D   :  r_t8 = 8'h56;
            8'h3E   :  r_t8 = 8'h6C;
            8'h3F   :  r_t8 = 8'h4D;
            8'h40   :  r_t8 = 8'h8B;
            8'h41   :  r_t8 = 8'hD;
            8'h42   :  r_t8 = 8'h9A;
            8'h43   :  r_t8 = 8'h66;
            8'h44   :  r_t8 = 8'hFB;
            8'h45   :  r_t8 = 8'hCC;
            8'h46   :  r_t8 = 8'hB0;
            8'h47   :  r_t8 = 8'h2D;
            8'h48   :  r_t8 = 8'h74;
            8'h49   :  r_t8 = 8'h12;
            8'h4A   :  r_t8 = 8'h2B;
            8'h4B   :  r_t8 = 8'h20;
            8'h4C   :  r_t8 = 8'hF0;
            8'h4D   :  r_t8 = 8'hB1;
            8'h4E   :  r_t8 = 8'h84;
            8'h4F   :  r_t8 = 8'h99;
            8'h50   :  r_t8 = 8'hDF;
            8'h51   :  r_t8 = 8'h4C;
            8'h52   :  r_t8 = 8'hCB;
            8'h53   :  r_t8 = 8'hC2;
            8'h54   :  r_t8 = 8'h34;
            8'h55   :  r_t8 = 8'h7E;
            8'h56   :  r_t8 = 8'h76;
            8'h57   :  r_t8 = 8'h5;
            8'h58   :  r_t8 = 8'h6D;
            8'h59   :  r_t8 = 8'hB7;
            8'h5A   :  r_t8 = 8'hA9;
            8'h5B   :  r_t8 = 8'h31;
            8'h5C   :  r_t8 = 8'hD1;
            8'h5D   :  r_t8 = 8'h17;
            8'h5E   :  r_t8 = 8'h4;
            8'h5F   :  r_t8 = 8'hD7;
            8'h60   :  r_t8 = 8'h14;
            8'h61   :  r_t8 = 8'h58;
            8'h62   :  r_t8 = 8'h3A;
            8'h63   :  r_t8 = 8'h61;
            8'h64   :  r_t8 = 8'hDE;
            8'h65   :  r_t8 = 8'h1B;
            8'h66   :  r_t8 = 8'h11;
            8'h67   :  r_t8 = 8'h1C;
            8'h68   :  r_t8 = 8'h32;
            8'h69   :  r_t8 = 8'hF;
            8'h6A   :  r_t8 = 8'h9C;
            8'h6B   :  r_t8 = 8'h16;
            8'h6C   :  r_t8 = 8'h53;
            8'h6D   :  r_t8 = 8'h18;
            8'h6E   :  r_t8 = 8'hF2;
            8'h6F   :  r_t8 = 8'h22;
            8'h70   :  r_t8 = 8'hFE;
            8'h71   :  r_t8 = 8'h44;
            8'h72   :  r_t8 = 8'hCF;
            8'h73   :  r_t8 = 8'hB2;
            8'h74   :  r_t8 = 8'hC3;
            8'h75   :  r_t8 = 8'hB5;
            8'h76   :  r_t8 = 8'h7A;
            8'h77   :  r_t8 = 8'h91;
            8'h78   :  r_t8 = 8'h24;
            8'h79   :  r_t8 = 8'h8;
            8'h7A   :  r_t8 = 8'hE8;
            8'h7B   :  r_t8 = 8'hA8;
            8'h7C   :  r_t8 = 8'h60;
            8'h7D   :  r_t8 = 8'hFC;
            8'h7E   :  r_t8 = 8'h69;
            8'h7F   :  r_t8 = 8'h50;
            8'h80   :  r_t8 = 8'hAA;
            8'h81   :  r_t8 = 8'hD0;
            8'h82   :  r_t8 = 8'hA0;
            8'h83   :  r_t8 = 8'h7D;
            8'h84   :  r_t8 = 8'hA1;
            8'h85   :  r_t8 = 8'h89;
            8'h86   :  r_t8 = 8'h62;
            8'h87   :  r_t8 = 8'h97;
            8'h88   :  r_t8 = 8'h54;
            8'h89   :  r_t8 = 8'h5B;
            8'h8A   :  r_t8 = 8'h1E;
            8'h8B   :  r_t8 = 8'h95;
            8'h8C   :  r_t8 = 8'hE0;
            8'h8D   :  r_t8 = 8'hFF;
            8'h8E   :  r_t8 = 8'h64;
            8'h8F   :  r_t8 = 8'hD2;
            8'h90   :  r_t8 = 8'h10;
            8'h91   :  r_t8 = 8'hC4;
            8'h92   :  r_t8 = 8'h0;
            8'h93   :  r_t8 = 8'h48;
            8'h94   :  r_t8 = 8'hA3;
            8'h95   :  r_t8 = 8'hF7;
            8'h96   :  r_t8 = 8'h75;
            8'h97   :  r_t8 = 8'hDB;
            8'h98   :  r_t8 = 8'h8A;
            8'h99   :  r_t8 = 8'h3;
            8'h9A   :  r_t8 = 8'hE6;
            8'h9B   :  r_t8 = 8'hDA;
            8'h9C   :  r_t8 = 8'h9;
            8'h9D   :  r_t8 = 8'h3F;
            8'h9E   :  r_t8 = 8'hDD;
            8'h9F   :  r_t8 = 8'h94;
            8'hA0   :  r_t8 = 8'h87;
            8'hA1   :  r_t8 = 8'h5C;
            8'hA2   :  r_t8 = 8'h83;
            8'hA3   :  r_t8 = 8'h2;
            8'hA4   :  r_t8 = 8'hCD;
            8'hA5   :  r_t8 = 8'h4A;
            8'hA6   :  r_t8 = 8'h90;
            8'hA7   :  r_t8 = 8'h33;
            8'hA8   :  r_t8 = 8'h73;
            8'hA9   :  r_t8 = 8'h67;
            8'hAA   :  r_t8 = 8'hF6;
            8'hAB   :  r_t8 = 8'hF3;
            8'hAC   :  r_t8 = 8'h9D;
            8'hAD   :  r_t8 = 8'h7F;
            8'hAE   :  r_t8 = 8'hBF;
            8'hAF   :  r_t8 = 8'hE2;
            8'hB0   :  r_t8 = 8'h52;
            8'hB1   :  r_t8 = 8'h9B;
            8'hB2   :  r_t8 = 8'hD8;
            8'hB3   :  r_t8 = 8'h26;
            8'hB4   :  r_t8 = 8'hC8;
            8'hB5   :  r_t8 = 8'h37;
            8'hB6   :  r_t8 = 8'hC6;
            8'hB7   :  r_t8 = 8'h3B;
            8'hB8   :  r_t8 = 8'h81;
            8'hB9   :  r_t8 = 8'h96;
            8'hBA   :  r_t8 = 8'h6F;
            8'hBB   :  r_t8 = 8'h4B;
            8'hBC   :  r_t8 = 8'h13;
            8'hBD   :  r_t8 = 8'hBE;
            8'hBE   :  r_t8 = 8'h63;
            8'hBF   :  r_t8 = 8'h2E;
            8'hC0   :  r_t8 = 8'hE9;
            8'hC1   :  r_t8 = 8'h79;
            8'hC2   :  r_t8 = 8'hA7;
            8'hC3   :  r_t8 = 8'h8C;
            8'hC4   :  r_t8 = 8'h9F;
            8'hC5   :  r_t8 = 8'h6E;
            8'hC6   :  r_t8 = 8'hBC;
            8'hC7   :  r_t8 = 8'h8E;
            8'hC8   :  r_t8 = 8'h29;
            8'hC9   :  r_t8 = 8'hF5;
            8'hCA   :  r_t8 = 8'hF9;
            8'hCB   :  r_t8 = 8'hB6;
            8'hCC   :  r_t8 = 8'h2F;
            8'hCD   :  r_t8 = 8'hFD;
            8'hCE   :  r_t8 = 8'hB4;
            8'hCF   :  r_t8 = 8'h59;
            8'hD0   :  r_t8 = 8'h78;
            8'hD1   :  r_t8 = 8'h98;
            8'hD2   :  r_t8 = 8'h6;
            8'hD3   :  r_t8 = 8'h6A;
            8'hD4   :  r_t8 = 8'hE7;
            8'hD5   :  r_t8 = 8'h46;
            8'hD6   :  r_t8 = 8'h71;
            8'hD7   :  r_t8 = 8'hBA;
            8'hD8   :  r_t8 = 8'hD4;
            8'hD9   :  r_t8 = 8'h25;
            8'hDA   :  r_t8 = 8'hAB;
            8'hDB   :  r_t8 = 8'h42;
            8'hDC   :  r_t8 = 8'h88;
            8'hDD   :  r_t8 = 8'hA2;
            8'hDE   :  r_t8 = 8'h8D;
            8'hDF   :  r_t8 = 8'hFA;
            8'hE0   :  r_t8 = 8'h72;
            8'hE1   :  r_t8 = 8'h7;
            8'hE2   :  r_t8 = 8'hB9;
            8'hE3   :  r_t8 = 8'h55;
            8'hE4   :  r_t8 = 8'hF8;
            8'hE5   :  r_t8 = 8'hEE;
            8'hE6   :  r_t8 = 8'hAC;
            8'hE7   :  r_t8 = 8'hA;
            8'hE8   :  r_t8 = 8'h36;
            8'hE9   :  r_t8 = 8'h49;
            8'hEA   :  r_t8 = 8'h2A;
            8'hEB   :  r_t8 = 8'h68;
            8'hEC   :  r_t8 = 8'h3C;
            8'hED   :  r_t8 = 8'h38;
            8'hEE   :  r_t8 = 8'hF1;
            8'hEF   :  r_t8 = 8'hA4;
            8'hF0   :  r_t8 = 8'h40;
            8'hF1   :  r_t8 = 8'h28;
            8'hF2   :  r_t8 = 8'hD3;
            8'hF3   :  r_t8 = 8'h7B;
            8'hF4   :  r_t8 = 8'hBB;
            8'hF5   :  r_t8 = 8'hC9;
            8'hF6   :  r_t8 = 8'h43;
            8'hF7   :  r_t8 = 8'hC1;
            8'hF8   :  r_t8 = 8'h15;
            8'hF9   :  r_t8 = 8'hE3;
            8'hFA   :  r_t8 = 8'hAD;
            8'hFB   :  r_t8 = 8'hF4;
            8'hFC   :  r_t8 = 8'h77;
            8'hFD   :  r_t8 = 8'hC7;
            8'hFE   :  r_t8 = 8'h80;
            8'hFF   :  r_t8 = 8'h9E;
        endcase
        end

    assign w_y1 = r_t1 ^ r_t3 ^ r_t4 ^ r_t6 ^ r_t7 ^ r_t8;
    assign w_y2 = r_t1 ^ r_t2 ^ r_t4 ^ r_t5 ^ r_t7 ^ r_t8;
    assign w_y3 = r_t1 ^ r_t2 ^ r_t3 ^ r_t5 ^ r_t6 ^ r_t8;
    assign w_y4 = r_t2 ^ r_t3 ^ r_t4 ^ r_t5 ^ r_t6 ^ r_t7;
    assign w_y5 = r_t1 ^ r_t2 ^ r_t6 ^ r_t7 ^ r_t8;
    assign w_y6 = r_t2 ^ r_t3 ^ r_t5 ^ r_t7 ^ r_t8;
    assign w_y7 = r_t3 ^ r_t4 ^ r_t5 ^ r_t6 ^ r_t8;
    assign w_y8 = r_t1 ^ r_t4 ^ r_t5 ^ r_t6 ^ r_t7;
              
    assign o_fout = {w_y1,w_y2,w_y3,w_y4,w_y5,w_y6,w_y7,w_y8};

    
    
    
endmodule
